`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
ZxTZQ0UsS9HXL+cye8KhDHq6JjsRKdBbt7/23hG3Xv4lTOl0WgHvvGUXhuq0kWEjqS5VCl4O7cYh
glsyN2zZsA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
D0MQ3ley4npGPCDj0uKNvxx120GglLBAwtK6OmuXlvAVN0AR4gZjPv9jfdRnj/KJCxgkNVaqUWhg
Egx0h1ObNRySsfchKqdWJxVp84ELTdz8SOdcwsqw3WYcma/EKO0xmVG+Dj5kh3SGzvvfDaBktFb4
bK3AFZY/+Kz6WaLMycE=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ib/FxVN0ZG+ayfRlBompcRYBpl17xB6BG0jS3s3PNdG6pBxEZq6Py/W4j+7qAMV4uf9WBeBuwU2q
HYo5rMUEYE6wZf9jBnW23+A53JEyx5cXbckxSK688vZaeemF9wCkbeVwfHM8QNbLc51/qzlRZboH
l7C4B2YP6+l44fhzNYY=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ws6JMsAbE3g94lwYREcMoC/8x4NmofYlfb9uHUEoOTvERSt6NSyR1yiG91nsEU3XfNhOQ7b/Wo+P
aa5UrHOplosBwW9O/BOPM9kStFRQfGsf8m20FxpwLUQdlNgNMPZvmEcAaEc+pN3iwPyX09CoU7cW
ox6RnElk1MI4OWVFf77mW8j6e1VlWO+Vc8LKoTynKGAP5hC4BYHQd27IInXzGdz1oVD4Bam4x0/H
sYLHZCISnOa94Q3CL6ay9xgNR41rtS98WTAttjEyFf8ILmaeESW6M4dGV3+EcdfBNzrTTc1nF75N
HxzYnCBLVG6X9yHlNRAwFRouHTyObDyWadNJzQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jKxqwTVbU6wQlQsyUl5EyNEaloyZKqOqnKP/oSoo8BbsW9jgw2GEmYOdPZbHNARjlp9P52Yzd3cJ
LczzuDU2cV2yn10WPFG38hLnucATA1ff0e8/mPzfxBEbAOPlzTkUFRukOc0zmo/tLK6cZvcaoRPu
DUI30FqzbS3M/o8XdN6yN2QOFivgXW0Xh8ycmXVtjktsm6ElnG31EW/2LkwLAyVftpL7G7j6nMnt
e+d+eKFIoGrxVI+7fida/LT0yaOYHWQh3rAG4GvE+2lORv2wy78727ZIirWNnQu8oy5qQcf7LAqd
e4MLtleFAxEV9eZP09SJZUSUNMj8waYaAU3w8A==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
w06/xQMdplxMd/DX9rImvuDEyUujJNZ5bclIgCUEQ3II7s7VZNfFQwqshU6852btDf1ThZcwb360
Io2jAnYs7UKM/nRMb56sYLBX4Y1+ufAYkpkHIcZcRICnnnvtYZ47grVBHrUfGA/xC7v/201YnNS0
c/L8l8Caa3RS8dR3ZckJnLnQOdimwEUdrhOFCxXNaVvcB1qFzyeB0qRxY/SqYktIcK0cf245rT6J
ycbkjnMIhAqvfqKdgoqIvgkkVe5grJuoukmw5uvFNcNJJ4EbH5xxoUZnl8pXhFueD3O6JeklVONo
/UZlkoZ7Ymk1otUl6y3wzaGnG8SCVGGtrmKfXQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 296032)
`protect data_block
/7nb8rrykROMwCEWAVvp/8ud0YPGcyoH6zTU/5zLnYpSsG/VdOTNZEJs90J8brUexS6Hao9iXy6L
Kzk2cSgJb0oSG4/59L2pnEmAzdaE7AkunMiGo+av9E+NI5XvJauPFV2YILl10T1gB3r7+9Gjx9TZ
miHrH9DL8cADihGkbi6eDefsbWuA8kHdqeyPtUgFfEg8wbZyVK34qlJD92iiD21Q8y+RF5EJTgKv
v8bsAJ1KfOCkNUMReFOzcbynfWr39L94+cs3kOtpN0eDJ+pjt+8RJ1fWG11zmMDR7UNgybOZAZfm
KEAletajBtEQaz4wfr2CYMXYcJm6ZSEG3xIsZDpVfCVM6e7A9wu7MBGeb79TRLgWr2YffHy5ZBs3
hASUSIZdBK5LCF3NyoqB3EtiTopmH537uV1unX/76PwoWO+w4lvxZUwtDZmqAYKQw1rey+kjAsa3
O1onDJIQEHwlX29iTexxNFxcxVbfwBIvKC9yXcuZRSLvdQr7NgEdrHlTVw3jd/zFYcr607r/jlHI
6BSLm6ttePhOauYC+qgK4tSZPfGIkD3xftZzfk0Hh+kL1zWKYZ+bZuS7HJHY9kTgqjfRWWwDYFVt
EFd6auVgxuRZCTVdrguWuzBF5uAmgscRZtA2B8spDaNeNBmW+RNyTNSmIpyrKlHDR6jZ9v+Qe7zJ
g57yNfvVgtzIe+yNuUEDVfIEDvcnVA4W5rMua0jBJN745GBDwEkp612SKjfAAJIhRgLSisc/z+gC
eSSolnkJI/4Zc1+BUN3PU1Uu3U92/evQaqQXdXHzR8+5bFxx61wF5nOdHD49BdFEOtQLrMwhcOF8
6scDskCLfD3leSYnTX/v5g4B0NUhDoPaTLyHjJf0S0s4/oI1n2ZSL3vYtvGuu4EkIT9N3BF7Ypn4
kVdeqTwXt8TKmgxSy147/nhllJEu3j3YJMJXIMa7IEjfRFEBt+kwCRkDoUZhGrlOKLd4xJfTpxhA
lP9oSSrH8SwPGFj2gwnNsNAlYrW0Gzq55e0e+BnmctKonohuulU6otF0wrB1vjqaesup00Qxag4O
oZ860x92NC2c9MC1wj8A8fE2kqwlbCAT6t9xtCIZI3cbKQ9rt29qg8optqaGqeh68AgCIC2Qqcgk
0+JW0KovdF/G4UKseXBVeHzWyMtCnIjQCfuu08gUnrgYxfUysoPdtd8hBUKKKXayvauP0F/ugXf4
wO9wI+K4jmGsPD1rbjnFbd1G3WENOmcmRDQIxaL+gSev+CBRa53oK3wUyeAA6RzPDB2YJhrM2kVA
KPwDIIoO3pxEz2YAx2Fu1S3+FDqm9D0Wd4gITMHYj2Q+/CrhcJztkiTTwV3AZaDeFUV3DXm1e27+
SqfdSa6TPoCTGTcU6xdfvTV7hlFufo2JN8iRMr0Yt2uoHo9WEGc88UrqnW7FV3U/dVmfdfA42N1Q
QEdjGl2Hllx4P7IC62plggo11MtcmgVynr5ssBG98hkuwCjs2aGRyjC5OPF0DSJgmG6ZZIW4CugM
/NJdzdr3Bg2XjMiriF39BBe2/ckbTv/raypQ4CFJ4FEJojTYAjg1efkUqy725HCv6muL6jdcG2rH
hPfE8v/ekamWiv+S9nLRwQjXsPk7Y5TEHs0O1qOPxnVcjn+cJdT7DyMWbXwkwDp85k2hj0aA4GWx
hWHD76rMqMHNu6bnaHrVTMe0JCHqNeMdq1aYKUdk/D56Hgn9ct/X1BWDt1T0nzvudJSTvtibdK1j
oDPxLj0DQDSQrdu8tqVfbR9Ugwzb+K6ercibTyyDYisbTuom8fVI3hf8cTOURxpFIX/zdqAB/cCZ
NmFZG6aQFuUkOEIj5E99UuN8teoa7ClNAI4L8nyrArjRQAPPAmHewD0k8hxZsYdNIxGw+y7lSbna
QwuCch+GpQ9OgoxosLYbqdpvgC0xqB26GNuxHCTgFeIecm+wQDqVGwZa2zWX3NPDPwymrZp7xRXn
d7O5ksRYu9hZU15jnYyIQa8qTvB+4Cpj2XrMVScCoVHNlk1uVI44Z1+g0D+JDkpMZIhoE57QXjp+
X+PPPmvhzeBqA1jh/IuOp1C63tYr5AaVuaahJ7OtAucVvKTKIju+qLJY5UVargqUTDjwfNKJ4pQC
r/ISqqhna42cqLyS/MP81qNvXXgc4ebBRo6SyS0PpmRPpp2h7G6YbeRA9uSONTwDiZKNZ7Wj9Th4
eU6Kv6U+9QU8JoV0tMqyjc31UAHHnAKpuviygVuM0PAZ3Yf0aXwkcR+7O+RbAwA5qNGK7puihOug
SzuYHhK+aBeOuYXCiK1zkfqHhHq0yRnVY7nM7xMT6ZntLiAQ4u1wRgMnoM1NBfpBGOdYwbtWu4b1
oTK/gwkXgbIFam1pZXXQ6Ne1F4vsG9U3OKFJd3OehyYRJBdeVlYl8CrWLG3w6sZUUdG3U/IJm3TY
SVLg50BSntUy45EAhQq+1wA2C9Sgjg0SidJ/Y0ZEdBYcfghv1sFEF+hLl8+ZhcHSxxNp4fyCI9Ud
7OsGFNnSmICT2COq9McTsgs0jOS4dKWfUZSWS32ItG3CRTNVwOdzLHj0d6QqQ/sOLK4r8N6qpYob
xZFG/heqCKRizqP4wgiMjnNnUrBJGIm30hEi4up/9JEjBJKGqsOqLR7uK505kZ37xmyxRerVtVIa
nSjBbq2XRaMnCIb0X0FETzQxo67+Xp56/tq4Qp6Bj3MJa39o0/sb7glppzlaV/dlZjoIXwvEOBMq
HMNa8mFIq9zYnBPV3/BvohiiFgcsN+kf++HDEHY3a1WGU6uddUV8kNPaf1bsjwQNgymcyXO2/tlP
Su9+v2ynmrydE9St9MBJ0LhvlXRyPP43Vwn/llNlaNgWWEx/Rn3uYL2D1uV+Fj/3he8lpXyxQGOh
9dVGAUJ96uOcdlr+OGUFuzIhnwCUw4QcLZoteA5Rn678CEMRyAnSIMA8J5qMpfqLqAsDjAi6ikDM
gx3SUtH/UAtLT1TZGYH8cdU4ybtmI9H99pEm+zVgstCdoSAgFYT/T58138SPxYANGW2s5M76rugB
/DBr9CZJ0Q1x/aPbmjg+sxmKpAqWrYDTIGHWcUOPP8QuMYR1RVQR+99dYB6h2d9lBk+HZUjedZO6
aJaNnnqYjyy9TzyhhS1nYws8iy3kqkF9t4oy8Fzo1SAVOr5xifjs54cKS8HXemQFX47clVmWsI4q
RUNKyAxhTipin+nvVjyaCUhmqDVf10kHXu0eKmwTOWK7pdpW6tKnLlcC4yiD0PtQWj7NysSfk+tO
4KpKZykZeNh7HX/PN1xtgP61VpZ/YVbq4crubMGGEp5LDuJh4ZN3ZLLOYKLzOVI6kRih07mEK9lp
r9UV0P85T4aZxc4Xk5ou77I/SlytTRj29dO4pwyP1Z6d6U4TAcA1drxO/c3KhQg0EYA89wCc4g5W
35k0adgACnrdJnG/+54sxbsphmnENwpgzWBmy2dBIeB7o1ZZ5PEL34dTm4BWCAxr0OaeDaxEHSHa
ElvjEwH/jgZX95anazDJoNV324U7ZHfdEQDoyJxSVwY8hcihNokOwYlnDNLJvnPINCkq5BOG+Q9s
e6ImzhAgTmasV+U1cw9iZGe/jbcTtOPN2S9B76QZR6a5kET7KJWKC2GBA2W7Rg7HcXeKBm6PGKMp
Wz9M4ZcUI2Bpfm5gyMPqFPIZw84WTINNuLNUVYt3K99bM9zXWejNULPOW3Gxi4Bnuh7vXva3mApM
iLsNCEJurcRYnXfZ408vHOWNMogFrgBUclbDxOC7n4ArUeVWbBBnkYTNeM0dtoFY6nLS1dizQXyR
KFt/QSoYmve9dlIr4oSMp6l3FS9J7+Tst5nhPVSwXPx3/R0sop8jwPwWCS9+YKfTDL0onDIW3sQG
xUqAi4PgF4AvlOk5Et3WsymKcWWIvsnvfhZPACtXI/q/raq145cj8el/1UgDsrhAuG3YlKcfU5TH
nuSSwpNlWHOlZBfmiRPsqMhlvuZo+HTUh0vRyvUrOdt4tsF1u6//IRbvhDGVstYq5zWlGd+vM//R
oOMotRJ9tqJQ5rZjL2WqbaZzac4vLwpWIPgj6LY7xxBddTx0Z1kAwKlnOIx+S5IEppInWPKo+DAq
Eiv/4HJtkSVXWXPAGVaYH4lLLthOdOAyBXQy01boVyDXC68G9auxHvrZRZqEZAJKrE0rckHvZmEE
q5k8G5ivfmS+ptoXlWScaancCemkLOQmkaJpbvSpSHDo/KQGAGFTMP9HiUQcE4LBic2KUlLQ2Ig+
d/aasLwX7dM8fyqQZdDLohBjP4z5dPyhWqGYaKXYVmY/IgaCKuKPwdsh5UbpUdRAdc+k+R6q8Eck
KjtO2b8AypnBhT7Jdve61g/QxNVaXk3/E7ylm974+nZVbPzKcYGw7dXrbhcHEIxsvrRAkZSVVFSv
Z8tErrhBY6WUT5qiAphjqyPCnieZkGONxFrMG3D9E+6qH/5+Q/QjVifbET3TsHTBl2G1Hkn4+/lt
jgEmqeAzeVd95NBzyuI1Shz8DoOjVKc7tSAMkS92Us175Acc1cpmOrr8OTdNUIG8tPaqCoBD9L/L
ej9VxmIeVeP4K6LHruI2uosO4DLrdqIC57+V5g1woSWEpbM0L6cAU42yWaQiUjfv53QN6bAh7iAf
KTEQONCGxFiKfFMgorZIrZs/TewCvyIJgr+k70CjfkhvB6b+9bJ0bT18ZdfbTORIy4e9z5ZPkHEz
kSD1h77w9xy4rntxLGGu0bZLBZ0cDtSoNpIUe5hzb+sh09OwyeXqH9S+kpcbuNajv4gkgXctvQPN
g7zkDKQCYc/a2BJtuxIawqIr6EojW142vJmNFeSlXr+LwkqqONE+Qei/BhTMBDyqT9ZUGiDNNXCt
P0Tkr/GSzJ9mG6hu8Jq4n1As0j8f05xCC0GhFjJzUUFUEZryzIwdtWg0hBocuL4O5cKri8if5xbU
PlrsNvFhz+DHhmlmDNIXSWEvE6ShAF0MdINSjaORtsdKDZ6Nu+FcpPGMa1cwc5VQq27IhFuoy/OG
SidyhnantqWYfc/ytkJGZc1kXRbRUWqfwktjzicmGXYcoC9K2C1vOTnbXQzMBwM4YRXpmYzPnVpV
iAUu3Xxt9mUblcr2CkPqytuD3pXros/7b+WKeanA8dg2l2V+mt8ie9v8cALJLgZHXICxn9plcMG7
XIGR3nIg/Y6wuOHlFlHdLwGfOuZlNhgIITsCQGGuZagwPhNuR2Xop/B9p82qmDDBwyBrcy6AFQv1
w9lAEcrlWkHylmQGZtV9FEawUC+i2gOquy6iT5+buyzDjCx8bLZtcvXEmdSFVXW5MBATVyjAGVM6
ADb+OWj7fBAu1Iz3WP879W0KlBCeX/ZlJmMWtFB2sc10lxrC7JnHkhkF0WP8Tlr3fG9yFsJx1gkw
u3H43yQvMnVzfGqOxPjNKSVVcZgnqWCWMdPZfiDCUZ039ro2fhpeRFjHCoGiUgFo0OSbrzFDtgq3
mtNo5v7NQOg1PElf9dOPZpoVOJVeNNIUd8LzmLMPVenR2KciEPJ7VYhutKgybkm4X5tQ5NPfCrHM
MaXlcudFbyJrO7BafJ1oqWUNSXd74NY7F/jpEIMSa+fkdfSUF1oI0vYwXbYWUgByBUsk9eSpnfhV
GQQCQmijqQsovewBeMyMJANoVGUHmHGkLB1j2Dnpr/7BQoYHdhfEN8eYO5Uz6COHL+7TV+qg4vvt
Wvuhp7zokF4yNSKDTgk1rIEpAU0bqgKxmvKKB/fwF+TmBiZN4xkFiwZ1mJr1wKWoD5CTcf0pDlI4
ImOhwlIu66Ubb+U1Xy42ZAb3WJZOCr0NI7O+ZYNv1J1un4TtqXkQd0UcsHll5crEAuA7f/9902Am
Pm29Zm134Wg9rmBWKfMuO0XIxJ0sYdX5OaO2dlyBlRaq6PxdARQzwm783/SwN+p4vQXg8PAzx+oP
T2zdqqNCeZQRXipqFtPAHpfl0z8ue6yppqfkLsje452kQDhDE2Uhlnq3kHCZvnBYJ7M/m9N9crAD
Y2Jz3ROK94i+SP83KldW/orbjwF4evh7KKZpovjTWW/XfyP/2ytbuVcb9HN+xAY/sQghSRHcqXyk
RcW1+paRUIPAnaMMaL1ur4upWvymzT5OCvUCglaBYq+wXH4iP0vcDcj447powqRVmEcr9VOPOPrc
DdseA1Yw+8iTpVWSi0+Iq3a/iRmWXIZks1CODkuaMqUnZRy6vcqMZ7771sElq5V072LUSNpcM8Pe
xRtIqgwFIm1LYHvgx4EebW+oUOVH0at2rGq1a+ee0cNtAOBSH5xI7T70w0IsR1zVgghCOSeNyaCJ
yNLL/CYG3SUG+bQJESRDWGhvHYwPgOl0QgzVonjn5U71v3y/n/rbjAU5HVBlH+9L1DKyuPrSKRRZ
xFUTGB7byqSnOk7PKavOIIUpnHenIqEi2DAYKYv4mclf/uwe937Fa/uxpWLGb/VYnME+u3FxiN94
JglCmwbw5LGAYM3hJ88brhPIGZCYJyPl0UopfeK1CpBTELmk3s0Db3108PkDeWd/92SxRKU38xBY
FNe/4tXkzlUn827TD5CbOhH6vgFSpuGNGdv9f4UWNXw5O6WcLDRZj8IYXTJeAVFuAd5k9zOKbfnA
wN+NDU1bdRbVirxdYiSX+O9oflQa8l9313gx0SwClWQUdocJwxwKPWPF05Dl/aeiFw8LIHuTAjVb
ctqS4HJRvs51CWpM0Z9Btifr/1M1PjM5/2mh2QQUstCpMHsGa1+O9R9czUUClZJs6STAueQgbcst
zJVgwCJsa3Tz4nj7JDldXxkWHR0htxkBYH/MkKaQRlJcQ0Y4wzi6B9dTYG9gXVP3kQYLsGOs3CeT
ULHEC7lXGIwhiZf0d5mJxw8fb2NkLTFS2vIPf9oSo/oam0uXtizhUuG4v2aV3s9lbYvXxiDLIAh0
Eoka4Aelzbsztn0+Y9ChAUiG7/7VW9GdQveOPquAV41WBFBCF3D73SLgnb4Slu2mf87meKZzUe3d
a6agHToRzmCaLfarQG8nzuHi+/MoHzJ4ok52LlDeHKa1TtgOgM8jOMwF2W9XkpLXZ79WH5VnWcV0
T1tglwB6/Fi3GE7MP0eA/rfqV2IMRGVE+QGFFJxV+mvTvLlHgLUJeqVhH2y3ZFl0dmTpa1q2Y8tg
ux5U5wYCm2lC3lurLXvXWvTPA/kLrKq0QaiJo/KDe9oDJ9/rGsIBkz55hHO/XEFAgI5od0VAvVbs
pMDhwfHUwBc9VCR1vDzR1ycYXNMY9Dya3RnJsQ5kQPwJ3c5EJtA2MW0gYu9kPofaWffsGvLLzr6f
lJYndzIkIinrthe/Nh8o7apV47jFTBcXpKOkPDGFSLNDs3SfXOlvrmJEHjpL3U1eodbEZKywc1Fy
pj+QwXj7SntkoA7pxFABvyVqQUDe0zDKNribLT3C80gPmzljjVP0kkrihB7wCBtO1TMU2m4q772l
K+Sn9c0cbthvMLcqFsMSXpNRNwcgDL8XMknX+Rgw3a6/q3rqKmA7F8wHU7OGBTDuYlcMpZsCjez6
fMr2ocrpDSajwsxiNTIrH4NTHBf5axDvfRsavpbQUEU1DR59hiMG96ctCDQe7UYSpXxuzhpbYH0A
1gXVrAmtI/qUefjekosctWshdufVukcmRzYwrzoG9hzJ/ZABoR9wTNbVSFkEM0G9I8NraoRbBQZJ
pcLGXZ5Z8obWiZ66+qcDmjwMUj9qg8rAP7I4dIDUE2q6t+TBvhDDiUx7OinH2fvGnH6FQ3bYd5sc
W7baQdKuvTDU7qcd6NdqetaOZyccNZW2kGmPgV3Oy6N7kid0HIjOrAQORfWW54dY9/CRLIh4b60c
ZbDI4fr7I3txuePWVCu5cIpnj1Z5zA5XawnkuEr56nU42namsBl7IQOH6NjRiJrcbWDkombwurpJ
2QgOvb0CfMprUpj5VHd5LO8A9AG4UuYj/3d0GaxWmRUskBdf8lUsQ+mJd4rIS6QocrzzZFeIoLrS
8/QqAn4aJqS4hrUx+uzZr+Uw4W/rgMjL5NPRwzbcMiDu+yGuJujcSKgBS4zKalQzMTQ9cqNtiwXl
ffmGLeDtNkbdH2rV0J4HcsTuUmR6F4AnkGOg+GlnPrmrheu/gJMV8LfES42e73fqRRxYOfe4Mu65
jT6IRiwJ/ixQXEsFn022hI03+3tTVrDbwpZifRLoQc6RGbV+xGZIM8RU87+9cfGclTokKu0249Dj
VwMMbcN3bxTECCSXIilR2fRwRLtrHTZvcjUWS15hkriGaqVpGEjokv9TqAPkFVgJ+6rsNpRz9v79
K8T1SEYDYtBMsoRtebUFgsuVzb2//xQ/xHJFubIMKODG4G26m4n3RONQslU5mGV1YQD8ah7bzhJ6
PbvVkVd/YvAQySq+KtiJ7/TeSHoCD+qOOyNG0dGF06ekP7g9Ab/jIfwNSZGaSKmYr9rHnzXzCgil
H1/6se7UX5UDV8wcaxeEwaJrtGpY6x7Zlb6FJzroLrOONka20Tv1qMNMMRJWOjy1pL4tnS2T17+D
G3iW4Qhr3nHsIhxnmHUwuYiDPWatW+8QI7Lj5m6Og0jVBwwDYHrjqIJ2BG9ayAb3izdYo3fRcGCe
TZmYJx3y3aqoMQ7QCrOKi9f2+DQUA6//9OqLOQ3QsVjz2RCWbp2UqMo0xp0EN6Y6DSqYIFAw73ZY
4XqN058t2aG2/K99RT8U6Hd3z0LuOfxuCklm/rjaWbU5ROFjWKLgODPSkINr4Pvb7HcwcZUrycxT
J2JfivsVnoqsx55U3/pBqW/bE4fxtuR0twcnlyC6BgCuYPT1i0RrSF2Hu0I4TtQ3W8bBE9kn5pk6
I62dLjfIu+4uM821dbuPrdsoohZf8sv8SC7IZEN4dT4Hayoulm6JWoilIH9zyGENf/eZfT2aH2JT
qaHwg+Xb1i0Yj9bHHMxTfJPFnhX6g4mEzlxgMFzO1IRkwZsB7oo2ivxtINScuJ2DsTjx6hCpoJnk
4cEWv+qk6LGvluH2quac7L84xsnKIzYayrxC3oH0yrrn6FX7Z1xJ9uAjZdKuPsoGFplQXqwTZhKk
FN+t+U3OkDI/l/zJO1a8ovpwjNYIDgPgvDhhCaU1yBCrZsfYl2/rIU6EMXL7oXaBaqsHL4KsgtAF
1WOtR1DVLQT7o07qb2LwtNrSCvUqzSGJAA1YGQvnkXvlOu69yzBF45UnyTeuw/Bu/dChWm6kMtjz
VEYFIUvvyEuFLsA6TjA861mieGfvqIr5sQGqVCG7UalSiz+6pzJI3WzpNw8hI+OT22Jq7at6kOve
IjRrbS3CYTNoCCtJA+rgKAfK4nOHpDanH9nvLQ5paycYJxwVM+8stZZBeEJ4OLN+OiGpgBZAWUuK
jYIiMh+l7Su+GyJD7KinsQtA/6n3+otsWuQvzmwZQ8fpZo3p44U24MbgxoVgAnQBZI7Azd/FI1Tx
BvvIeSYNxJruiBuEqPORP4qERLcXhMX+gH5el4YE7CuO3AUIonIs+vC6z8GZExgB22FBWG68wWov
Lkxro0wDKYxlDSIL8h2VM7H5mJnakmnpWhHVYSnkWzgK/AkssbJNfOsat7kb0PEzeHTcxC1irzxC
+WL68BW3ZzQyyoFkRYYl3k+Ucrlrp960uE5PBHsLG9s+WMM8w1ZjdNdX4a+GXcX3YqMmsnNUJJ9Z
QhsaarasEozpwqHlSxxK+kihPamY6zCnwADY9+KsRKu76pZ6ioSe9A/OvV241HezchNVcf4Kb/ue
IFjpSxdD6DE2nn5Gj62GLO4ovk/Un93+aptaoD3QBWfZxA8Nsyyc6gkcTvk7V5xrkOyVgYbqX1ds
Txd44m4ASAzu0SyqzQ84O2eghZuwl1e4KhZwnaKFvXj1FSPsphJFpjEpy7ECUpyt0XGGlFKysoHP
YhRdkX1u484YOxz+2/0WW/KhGXXAukrGKx96xdEFCU60s9eiLtuw5oK7z0ueUU2KVZTE7TRqoRtT
MMKf01khEOsS/2A66+oFrePPw1gXcngFIhJgqeOAimm93e/V2BUqQmDEB1mQjFsjmWXIRwU3mk1W
Jy5R5koG3UKCD8B+PLbHIzkaxQlhc54fpH9+PbWTIRyWeswKKbeOvM5i+IUlapdMCEm7ohykjp0W
ST03zVA31u897B1cKH1NKaf/lm9WluuvG/wNEyHhEsaLiGM8Vn7qmUBAy31++8mHvcCJLCNzs8RU
P2PDsHaRnyzGgc/ZLpAaFD/vj6BPI2uFka9uD0OJ2Odbllmn00J4V0hQoFCxjGqoT9SWrH92rc/u
c5GZj5TjacapzRggYatovU8pz5xQnDjLOIt7ktfLThsNmV9E3zikQNOKDJ4HHDAAarY7DG/11k7k
wzg78/I6ZxmWbj1We1GtDkF5j/FQHEAkjgYOrYD5UwnHlhUkOdDnMJch6+PgolktfN4hFvEN1LCn
MvvUMSfbisPJXCU+thRCfor5ITKvEOVu/iusfihFOYjj3w+PK7lhpTcdXbxlOmy/kPPCFvAUkpyg
/DA5n6jv0BiZJ07vfOLo/1XyA/f0Ai4DBGaHyO2xgfFRA/b39cqD8+9cGnxtUoV+ito3WvIAFA6n
dLozawRz1Il0U9njFIB2gyrCyorLaL4PKnuqzgPX0jTUgCj2ufmIYHNMVDy3ClWHN/M/xDtv70Me
2CndfltcAYffccpGZpsy7tKmLSkMlFWswPOx6qtUXw0pmM/8Wze0bGPh9fPQpoMWFx6PUTPYzdIV
XOSg4wKzHreVmEzJwezrx2GOqt3mqrHKhXYlIswcXGVaedrwTr2rkneTMAFk77ev7azUT14QdBOI
2PII9X92O3MCdceKAJHzRkTeDPPLRjdClMdKY4Sn6oL3eWQnyw4fkeA9JSnuKEAEkyA+Y4TA/K+5
fO5PWRv8YxtKkiy54wdI38lmlxAp8MD+YJr4DwBzypGgWSy5XoUDW1qMKyhPd477rdsxxh90RHZa
OLHoriE0th4GZ6+o4W3XqCcKtVAVBacUBBWnj8c6S1vSHL1g4ksmTr3QCJukPBt55xEifLquKE5p
pKuHGi9RRDMVkVX00T7PDMhkgjwP5cBYduHZVzfGPVb6za7FpPx53QZOWramAabCM2DbXIl7wSL9
dhYCxfL9eUB7oYd3ZvWQGS98fdo9XVubrbBOxW6pDfe3UnPHlK9UtxYZJ/5Yts09+OvCl8dCjgth
PAO9SfbsH355Cn3QA6AY4MJgvFSU4HZoaDsPejm6kvn6e61AP3sKznuPbHtR4VgkpO5TxNDg2dQ0
gxbNxJbJUo/yPwUCKdv+XetmslM5Fp47O1fcXPsxmrHNeujalpo7EI5SgOAnxUDmyO4TlKw+uSQj
1kDNia9u0O5TmkPiGO4SKCqzmwZRozmoCOfpDq9bjiClr+gaI+6s/feIS43z87vWVtebfpTo6LEV
YkFc+gLVRAqVkaBLwZG4gE9vuEgGNSkYyXTlANxIFP8BLhq6Hd+FoJkt8H2bNOmrVCKdZ6PGSqsU
O0NFFQe31qXmer+MIdBj462qXvrc5SHMmF51J61P7gxHcDpfiUEMMLN46/lEfcaVEDh36bNwWNHJ
Bxh2Hhst5jmZ5GY7bonlZXYe3714+1fx2kmlY1iy/eKCltYz2rU9TYpuUP4BUXBNFf7RLTi/WBmX
w+WHirhXx5IBpKBbTLlgOUZLOtvc/o8PdRO5MMojILnVv3UV6wuvTrVEo2ArGitjIiSTYC5851LL
5N1ACk6CJkl8aRGssAM+3wJkoMXgh7tzM8l6TYwYUCAj4gWorQmsT4e00l0Rf0fg1DaISJFFOh4w
eIJxilQ1wuvMPmE8FwG/KUetL2k3/E8Ivy/F1+agR/NtTrkX5l5Y9dOjf6CO8Hkc2lQqHBdQKYzv
/9cCGd7SFjWJ7I1S6a69gM0dDWHdXDK/+LvydlgG38b8O6S1rUOh2GN3dY41JrRmyKFWcqle4r+y
fuzaGh14g8ENJ4jrOKwC6cn8VVuhJ2DnezyZavt3jQRi/fRUcU9ACj/ZqQoMJyoHPmzwgPnJAlPu
HHC09F2d+BIOQaPUgLMGLdsXH+WH56REFfgbqX9UoOuvLcOkFlExKvrGlf07sYqGlN+1R6p83UmA
/FiC9+YEf8koydQ64ASfGN+czR6aD3dUaM0CJwT2mNZqx1Vry9WueClbDLJZikS2/AuSs/48qrNo
CnP5cq90pT885+Yxb2oSttGyIKEfHQn69lONX5VhckqFQRZW6r1MozYnXYhEbgTC5vnzdTlWlkRj
LxvIQPswr5eO2bUBuVEPg0dYUeer7/EL1mZj771/T793YnghqWBeyube8QSS68hfwzS6WOz279XC
RhTMHjC+pYukZIG+u/pb1oghlZJloOyhCegYvGm40F+CsHMgmU7yQbsMeakMWi9+CY/PGE+YflEc
i6I7rcua3DtyGCKURtnJzRvRkJ/h+NLiCx8dNFZD/GjcNjiZ2OTYv/P2fOutjWD8TvBjkHG3DuN5
amPZBpJIkLR3S33J4REi786i9i1a9d0fn5R/5IEGTuGOpzi7jddDiMOHSWBP7l6zqINgdFjQGC8Z
4AguFsHXdbh5dSfEt6OPohnJ1PTSvHcGzCXweplS5iPdfrwElR057m4P0cxTh3wZaSDe1Daondbj
KomrvJTKisx2XePPSJ6jMIivuIwXFjPo1WRqYiwFPU69VEtvgcQgygGx1h4Sy4bQnAgnvjkYBMqY
LuVMwWTZ4MPGEtQoayGhh+fMdBKZzAoqPMjEwVfsZNAyAr9+dIqlZcr+GvsGRQq0WFUCadYyv2uG
co0ZExAHodI3D5yWE3iiTVKQ7fe9sKw85OTPAOl6ztM2AUs8AAlHw7nSSobTkimDWiNY5lrFf7Cq
J28PDrB36XzQCOrKqO5mXPiadvGWDmq8GHI+cTbQSSQ0Q/ASra3IQhbxmMoeM0hq8OzF+Pf7BDDL
gM6g+/sxdMYHYNEHmP2KiZ/cgprwBJO4hnRd8MFFQFSP9ZGxZa5/Od2f+D52Kl1Cn8WrYjLCjfqm
tR6JIjqm+A5qILQZcMHElk3J32NfNq2yr1BTJKt0yY/kVMZ/exEFbUp41sooq2ItqRY56JiL74M7
yMgqstsy3xLhIX7qb5H6bcq7OyAmwh9Dbp2DR9ZpzdU1ezR0qIBYPhZytJLL2ozgMsVNq9SLO37y
Xur9B+xwYfiMK2ezv9XxijpU8/7i4GuZ2diYk/rtTkck0H+eAwU7yWQXVstXKUSBmogM8Duxcnje
x9eS4c36ucj6j+aS9AmT4ZtFjUrmkx4uLCo4uJSvSZ+bdPTQsIbLihUM0IefLccSJqbLFsQQCrxo
y3Sqb0ubM1BEGq9usrvEjMm/nvrYM7Ve1YXxLt94eVjIPOdE39gwc/ICPnzTF20sQi9kYC32Gon1
qKREe/P0tlk4JrhZYpMozSrEZyhoG2RDYe4YGlpvjKx4HNlqxQdMox93EqDNAWFLEGq93l8GJW/s
+gibnpJO9500odfic3hiP/W1bddYYrWWDwc4InJxiIeFPLUygze/zcQ92cHRBgeHN2NOaF/gfgtY
IXv8rJ+q5DY87ESyQw16x1N0MUHl6fwb+h37wi/12iOgH7ZkIG/PqrDX4jzef5HLjEaM8sqBU90k
OEPl836xNzKq4HkIolsBzAyreB5ULi+Xq3XLm+FqXYXPIHTKABMYbR2IF5MoTwaI7WjmcQSIEElj
vsaqn3LmVFf4ggCI7Mp6sBR7el+eB8p+FWR/ktqj2hNTltrkZgQCw28NJ1OThpX1LyYKYIS92Z/q
6lcemEF2TaVxcnuc+xOT1/7geLLlJeyYeipr0r9BE5VyJL8VNfvYtIKZfPU6AVutq/e7Z1t0nxc0
+qqSolb1oJ4RFhJIUtAY+sU023mJilLZPaAqvikYw5vrRtNul0W5voUO3j5aJVyEypMpD4hgASFc
m0BtvAHdO73uwr0n0rHZ0UZphEqjv0wRst0w4koxaxOY1puiFnW7xP0pi6nRq4DSvZnAEQbzFzwJ
nFjgae/iS6RagsrwVSTukBiHSjzjUfo9rwJmpeAtYd4MahxdIfEIAVJyKoEoZ1cNYE5YdSdMDcjg
5/GgnbZBDkgpL4mklugttEh/6tWSF7CWpHpk4/BMoFbFnj9S6bSOa8x1sALejQbl6A395e/nMX9+
oGMmhyutCdGek0W5A0M8PKcTY3Z0rU2255KjGCyNMA1H4ZwYeKretc+6A1OA6wAMDEz+wSjM575W
OYSq+/AY2iw4UpT+02dbmglLLSeud9hBCqLQ4dyJdS27dxq/yz2XrR5vhqSHPz61QqdWL0SfjIzL
XrTwQ1H6BanBXUVKWPNEqW6tU2/DD9tMrPBqfzXssjmDrThWIBs2tiWkToP8JzPfQxXEU+uqh7MJ
aqW2lmBDSNviz2lYbKjXaUytAGyb+tKwUJKDcfdA1xy8LHi6r3SqjMJkkjfYQT12M9+Jd41lmOH0
sVtO6Veus8cN3hawR+wQiSrRZGzldbwUH898LvDyKoLufwqhsbOBVtSgluM6tnUv4P2YxoQx0gCc
szDuzll1mAqRJ9i+Rfg56/5jyPlHhIvW+znqmzf/B9Vw1nTZLBi24tHcUn7W/1E8FAsQZTEKzptt
2tN/jnjNNaAh1LfYFl71zlE6GPYdap5qB9ayCpHK/y81If62ROT+qLc9I5QNpHkqNWJbRsWpKwwL
4qMHZ8t4PJeG8ZOo49hbbe8lK5s1wDrLmOs28T0MhSjamQmV8SiMjnMzK032UYqg6vSxlHgMxEyO
4CtwFfxkEG19WBz/3CULnjgai0LBx4RziXYREBCYG6/PJezvB5V9ivB34SV+D9c8qezeJ8vmiuol
vv8AqmrCzWS9uaWmGIKa0AdC89T5s4SDoFm7NBpgjdiLpISPCzVtROadOnHwbJxEZ8aspGkHetnJ
cJ8yCgu/cnMA+8rf8DmxdBcdOG6ZbKoeV7KpvD8RhNWmsQ4O1AN5YUUzXmBKXX0TVskbTVg/9p0t
WkWOdqvB7TTSBBQYZmFcx+oiwXDVNag9by3yFnGV1UZmfe7xQ+AT4Uy1gmYTL3+95Qcg8e4Xjw9Y
5ChyKrQzomwx+UPxD1YRDIAlGbC1OAoeBVjGvv2CEdqJU2aCYhVVeSXsfOl05ZWQrhvngraNxF9A
8Y5yGARDk3QNmBdmKo0+TImgz4w2Gfalllvd7m4lnhPwqE1FoGlrsoDhDT6MhSlEL/i1cUDV6gdo
k7sm6a/BoaK5y/PnfAjRij+cQbNA3D/NCRMZ2vo5Qohziv+mLgTTr1m2o4Wwcc+dZ+fDL0rwAy4k
GQ2pR8BZ7WlrpXbTZnVT9mwKGbzj9z2XH3GpG3c+0R/ncmoLo3+R+lbI+rZbmpVT+SxFbSKC4urb
PiRgavP2iR1pPT3GMdCIDC63hkbGkT/iS8vbtrUUDCDOTOABhLhHoxnLs5R2BrIb6iN5l87jm6tU
enF1ascRF+ZRoq9fepaxOHv6OIBFPSj0mcgzeyrkpMBvkS4V6tNTUbtShftOiHsvUHfmX+7Wyew7
bnYCzr0W/iy6WEJDf+BUtipw6C1CH6mr9yWgCV2u3Whr45+YuEsD5B57SDUxOGDFVrooapRKCfuZ
cfAUxlxC6hq/dAeckzHywU1AqW9yqUnRJps/5qESyuXE+gPBFUPh16ciwrPylJRvbdjbAlF+oDP2
vkybmudGrB4EQXDwHfHEupe1Qh9ABKcqHmBLjFvmUyRnz9wOPotdig9lNeNSGyjWhAJHxvm3+RvO
/adlsRXRNSPcnBQLiyceYvTHabLdX5kHczxrgo69Ek90xcpuqIttAu4xkEjsc9EEmGcrUrtq6arL
ax0GEa6CU8plBHtpLA6Im6Gnj3/ec+UOLUWRXoQz+VaavIv+qfI4QqkwO5bcw+R/5zyqXsaE0yMK
BzQ9aJ4/VXsVhp94AKuYWEAIjDMO9TXCro+HSD2MKUVW+6g6mmPcAe6T2s9vwA6MRI0ut6er9rxW
9gf0k6U2sHrfFpohXZ2HlJfaruJkcQ8ZAy0rEyXVw1PkLuBRxG8dnHQubQl4d0cyjYkwzs0NzTT1
Xp9Y1aej4diQxM/bMzaeEOPYYNekzhf+DekZLEHIJOEBqRdsFHqJQaLJ+U/joka9Cr8U+mJAbhVD
cLOROfQzkis7+orbq1pf/ovhiOkq8DoRFu72x/3i6Fndoc1Uqfo+UXIuQEYUbXyEQdFX9/n4zLX0
pBXNKSXx4hFeArIBz/Gj3MP6y6Y/IFAmhyJ74L+pTq0qsM85K3gyaYFXalhTwDuGGdYGSkHwCsGb
HVQBShH0GlA0ecg9e7RL6DiOP56Rl3LTo+LLXBtlHMZguiTMkSkGwGaO4tZJhlHo8Yhqaad5RSpD
0U1Y/xrwdbvJQifItsaPvacI6oszTgrQdUUuCzDzC3mjr1BSbL5e920b32pz4giBUKtr68OUiOD2
LiWcYpa2QNE0mManj1pWhuc6xe2egOTLc/PY4iRTLvqO+aQ/7Amw7qT+w/IdVa2zcGjSfdqXfXrO
iU+/OXEmvr631eSsfcl/sKmQRxHL4Co1isBrl3aSSJBE4Cv60FKmf5lRzETl95t1IeAIRcadjAMt
6OUwkPNrzttGnIFULJkaPhvpkvuZYHS+t/Yai/ZIO5fbl8ZuI5vhd1+uB+Jk4fR3MK9YrWGYIXfU
lsB8wxxOby9NrrX3kPv9n81JX5BvJac6piyxmNNH2iAIQvvidMDCms69ese5vTIE9aGDqeH8Sj+O
IoA1KMlBXMZapBSuRFO2ecc6wwMYjiyIXsjm444bDKG2ZlNthW5skg2EJRvXSkp1ZQlhv6wLOcos
nnwZ/q4zux22+VFg5kqUC+zUipeb5DvhnZggYZmCdaPBqLM0dYcHPqwd9Q5PI8jKDnkIY9iJXsCP
9A4Bs1UHtkxelqE+VmFE8xohc0PXYpXQKyRRFJeApFhCo0UMDgQGJxCVcUPmgMhJNww48PkJFCR0
NFGVd1ikVATrmBOSVLkHHeeeTkSlKvQWU0lALARIpZGRUsroNhO3ymdUDD2WSLVEBsTjo6/dScva
Z/TH3OloMQl9rvo/KA8jIomViBLGT2qxfx3/F78wTU9OpaEXVjHNLT3MZTWSLsiAlxaiUI62VrQb
Wr8WdV3zJaF9/UWMDZcXnrx7zUWAmbLi8u3uhSB2CArKdzqIZnLbwaowbbBUlf7/ZLVl/xO0jHQM
kXNOHIfsYJFjC/M18kHB/dATdTLG3vJCsoksT8FSJUmc1shyKfH6xw2r1+a/dxYyHPOL7JlBbPz+
enSFsX0obgm1m4H7RmYoGcffPPMsDh5YCAeXm24JmrTKVu5PVpAg/WLYvLRUPnA4JRXnn0U0SpjT
vHGHtlSzZT3sBHjws5VB95PTgxL8IeDL3ZEEUhbw8fSoK/HFcEp0I+eLKZv/NfDEPJ0RVUvrJDiQ
7M/Bslcdo9pfQDWKcPQs5E7p62T45cpfvDMpL3A3nMzX4d291Cre4JdyOuHEeR0p9Zu6VevXVyxC
BNZq3sOAr2F0mlwnbxFK9+UxN3/yTz2ilB+oKUbdTNjBKnlAb1jAvMgLlixy4sr5/q0T4xvpRXpm
ItKfP3vgsHogJATZgXweE5Q0W5d3rm8YmeLCH6p9BwUhFmJZ9WvKkrISKwJYDAl6HIHFkFgjkCwb
q3cQMmAYSqyglK2VjkBOw01C6cWsLqDLPuRTeWDN+5g60b57ealAqX2T5NVNoqrmFo7tdcO4h2Nz
VnkZL/FIB1C3qaBMbXMSt1Uu5IS2IhM8ZyZAPHCGl7Fp4hJIb5SphhnTGeN0lyIh9V5AFFy9LLgj
UexQtOgRZCaZdLLQD952tXVyrvi4pRXam5yc6DH2AuObfdbGuUkeEVnYCa8uF2fuJ6r37ZeWDnEC
/iIbX/euy+uWkRN6ZcFmyCpquiZ9lSXP5beFwTPNQuPAMHx37tX7INKmONZB2eK8sjV9Gk+lh5DH
tzekdtVEHd6hgJsiWpARHHtueA8NteVSAodpuwKLKWthSI2usvxNhXewGdKBx16DQwoJ4G/e+9tI
yKTKA6m+IrXcdCYj3kjy6IjEQgizItMSzy/XtcDUi93hUTKsCrVC4me9anMGjGcvf2lBtNDKdQtW
iiTZnB/m0fghrznZOQ/yobQlgo1LaSQ8SVZMqERZg7UGeUwlpolY8uVMcUHqlXw9qBbj32mZ4rVt
j5HGlH3Ia12dDkJ9Qp+LIL3MFVnKLNmso2U2Biy9QzsUzYmSbiY5kizZThLl9Ac9voVsTi2Gmufu
0YTL+yXiwyoDf23T/+vuYa/trp65lFxOByxPf+BBO45u+1zvLATjj+phfeVQeMmv3s/GQmr6veW3
XmmUXBLNmLMhFKlzLx4hw25o1Sbk8vyHNwJStQ2lPcUiLc2hbQG9K1SLDaYLqMjx+ziBGlMbqyMu
pZW9jJzClsKS9b5lZqUPy02hqHUSRpkv0AtwtGjcqzM24I5n/v/qTkF2YPXWXpAYkHDrAV6eLv57
u2XByX3PkWNDXHeOzQTdAFzYpKDvlez+ltXXBqEIUHrClInYjPT90j+IW75yDgInoJaSn/SQyICX
KnIFxGSH5Nud52nWbcWYeA5I26BFVa2nhnNbz9V7mBoDQNKNbOzwcNLJJYgkz7yl7ZYc5E6m5Cf9
pzzfkTIBBs1UsUTTA8dH0dikPSIE5g7IvLG369x5IDTRPvIF1LOQCGGavsyKUYeFCHY9ul0gkBGu
YCDEqM3EHiVyw7ImTLRXbfrfBxJyA0d5T2e50xQ3FrM0t6WR0cJCpwlfqi/XDQyLFhrGjG+7APk2
acFmKZ1MlzW4m24RnckmPfxe+z5thNOCUMnztVOsgRbL34z0184sY0nvJAWUazG1n1a8mza5tPTw
mwGje2NcfPh1P8vj9y2XuGvXOaB4KJPEzbAG8zuQ9I/LJxnjozRSMMxiuZw+nr3P+H4aaQdLmCY/
hsgNHI+A47Iv5kt4mAFGY5P7YJXQdKLE4Y2FWkobEdWZV/jk2jKDs+YFPtuKydy9vi6SrVuX90ub
0XiRaOWof3IRJKGWEvc9z2FYaO6wMWEZ3XCaPkxeFONhzJn5Z/a1M4bQ02cylHhxtZgbYYpNlx72
WGJLyflSD2VxHAlMcuEOaMuNU2fcgLbv3t29WEjAl8UGAA/I4LKhO7FVfVdk4C+Z7uqWiHL4CFNk
pfRuoD/fv2USd9eK1jsRzatB4exyMcseqkvgNT4OQuzMVZAkMFiHKOHiqMKnrYbRSjaxeMrVDDEP
BChj4KnOQNXcPaYDm+dqJHrCa5mUpa2JVAsqg/MCtczoH+WWGzgdvtyLtupDAp66/Y0yg/GRudTX
sY1EMC7yCpRtSnlEKHO0qfTPd728UZrBaKN7+g0RNXQw4TeB+0CnwCB2UD1x7344tTH+fIygD1qx
IXA1YomZUIwJWWrzI38JPJkiK8nqEAUvgD1f9Z1MYWG0Y4icFoEBE+5TTkO4HpUm7F+iYhOJ+ZWK
ruUdsIh29BmlDkS031M57sLu2XkLkRNp5QoGpx51nu8zmpy/w7z784O9ltR3YAkDhcDTOjBGvTlG
tJbdx9uk/5ztmgeq00KHB0OWgp1M/kM8BqrlXLXdERyLrwejsCjyxCeYdN+9TnqReN0z/2mYBV1o
qjtC9N/9EMFj0frSM3C/1PbXlz6s8hkrv3GZ+/r3T6uwx6cXh0EsJMhcPOQNfZ2uFa0yoQ1IHGMr
9Trs6IdwiJI9bZEU4AEyGicyVbYFE4rWCnvlR2xzev/uD/eos5QHNWskJUyHAKT54BwH6UljbrJI
r2A/WjKt+HmvKDVGNBVjpW19IS1k0Fuf+tlTXoMhB6fE1amE9u3xif4RLOJiZfFjq8IX2vkdu0Fj
6DdHnow2h9r32DE2f5yzcC35y/vDwp0GY52h4/3h4ihHG46nO7QkobCxY04zJ6ygUv4w+vPN39tY
xbmHIxGsy4qFy9ec1PbafgMg5avIm8wT5RTySPwFx+MQ0+BPpxpHrAVidxbW5zrpLOkpaXRzUsVL
jay6x3jnNlMrO+OrVfDWQvHCMkFPEfXHHb/4FfAEWlcJL26ecGO+0QDzLYNO+WB9wl/nDP/LVV4T
f+0F5Nch6Qe6SPAbNpmYxuLNxdtFQUaJmlyqoNFTeFnRi+A3OGdmivjfXl0ODzhLuPNOKU2Z7LgQ
FNOX9znzeFbKhv+QTyoh2JqZIZopd0Nq101PzbpekgKqn4rinLn3FJBvkJQky0pRB/Q7nNCdo6TJ
WRq+YtrZoE8CvhZvXrvaCF1tnjWtup9IOWpZUBJWVxTAyHMdSa5AhEzEufBRe0exsbCfAeGTY+7b
gWsw9yYw8UzMXHQUP2gvseXjLnMWcyrsx8RU0pYEplpLJfDQ1D0zaglnA+d5/Sh9YyKy4S5OlOeS
f3Q/Y5F9FKFAUh7Gu3vnqm9DMRGlnqwCVyLKL/pnUU1AAH9/nBroA7abG3EKi0+3ymt+qOuT49D8
+5YOj6fw5iPvI+ANhcLd8bUhGLHktm/tP31a1dOzwuwL0qbrOp8Pa/4iqt/S05Y1Hyi9SOBjbJoa
DaBpuY9jZCSOUWiQZoW4lywGnO0c9eCpNHyZ/3XZcTbvAqWY8wK+DXjZjan7w7qk7aK4UDlcev9Y
lalqYTsz3meSuJ9xJyGASZBg952G9UalhNcV8rmQDW5fpkz2nl8Yjv+7408757zZU2BgaC+40Oy3
+j/SJNPwyANUM5O3GBvxGs+XaJicFE2AWbpOhvGIO9MRi7aF43LUBjIYhH01asKOHAP2pHNXDKZI
9tYWk91HKdS6JYK0SWlNSiebOve57ElYP/aKfQ3BLg65O2WwEPBb5R2KhovaT5WNLAs4RH8QRiZ5
2UPDrrFcXpp0srurRuN7r/HxA9KgZHWmir3hkvQL8+vqCzLmjQzT4ohBKj8BzLn7KoBh1gqt1jA0
IkZyfM6iT0ixxtCnmCkpCRMk4GGRbhrj0KbDu/GHkwprmWxD5Ck8dWiOQ2vC0OXYKVtW0Pqk1BIW
z5TX5EIHSH/si3bm8SUiQbEgGDvMjgCTStNG3OSipjzHf48Uv2ft0qUgoAKpta1eWdHZK9hscefc
XeUceyJYmD7zSAR3ps7HnNYAQXImi+eWQxGbNa1Hk0EqpVzChuO5gS2KubERzIK5tE8YsrhqPFwF
8cF+k18MJeJICtkIXtHvGrnNvad9NA0Wq1aN1tuBnc3l02tU04SkILqq3dmzbKxi0YuCvHjAymVY
c0YfWwRwQY/N5m7HjHPQwdngM4hAynhQHltl6h6uzNZSYb26tHgypJhVGKJbBrfCB685HS6aVuH7
T6v/1HfbwsbTNNID4ltGtKHsih7tGDTg6ip32B9+1djZn59KYhvtxcTN8lg6OAv/efrW8v5TzXFA
UsWoXwsZoPWCJlosNZl4jYGQJj4J7e0uFJ0izV/2N9DMKsR7fYikOV3Cf3fdmNkjMSp27LW1a/RA
pSVWpd+2xS40CdY8cTSpiaadc0BPWyMlBThascHjb0oVttcAnxwnwXPNAKSkE5OyV26ga+pSmsQD
tBXkGsVwq3tbJ4YVz+7eYocFvNPbijxWmwXpsmHlS69hk8PZaOpbkf+olNkVN0azIwbXR7p1Vz5K
yp9yZNVmazLeSIrHcMMqyT9BpO2PqA5S/qwdqwdcYJDkz9F6xvsw+jXRjreEQqj4R5gx+oXnGVLI
oHpPKhfEr2g7Mj1yRqMBTcDXpaZj5KBcZqdkKJSs2GLhv7pFOBHVmSI+by/Zs1QIuL8chNmnfnNp
d8FyXZBm2PTCGAXPpUxda0NHs9Jx2W/mLwzHlLcXQ55h+3kR1qxjVXQ55vCooX9JX+HPWuzon9+l
6t+5i7RYQEogtWL6O9MV4IUMaFWgBLC+g4uV9+tjUFRBwaefZuWtyglpeZRBKcyqAv3NxiXJ3oE8
/2B9WyTVsRcyZaYCVheLgthEJuVbRe78cv08jpk56g6n3r39OrODAgay0aPJufDFca6VChvFS5/D
sKIzkjZF+xOSy1KlGhML41S+2o1+2XtALOzWCUQA0XQ+9wfHb5d2zl8L81uITsCgrujT/PfkDaTm
Lx7CK681Fignt/PuEGHtfV/lmHVwIzuvW1gx1lvktksTq1/q2GbPkxqPudzkIHwZ1Ik3vKnsvVzS
ATrNpGFsEMI+Wo+kzIXnnpIF3ax9AO3B48GqPGJSRHBET6v4rbV6uZoZOxxHF4n7HoVBPruaYpoG
0IQ4qI6mUUNl/SIVldBdDgbXIst+JdbdYQ9RdgiEmBNjXn+UPyQIDjCmcvytcVovxAjD9bW7H1mn
QeTVylLKUqeL3gyQpNZg5X0cvw/apJdsmlW5zRBmsh54uvcE7s6wzrjFpkW4g/ZBc2wnYYtANxw/
2SrQSoUoHt+6uhG0uFHxzTV4EnTBRtxmFwx+HgLYxqZ7Dh5H2Q8lO9JJdzo1aaQfSIsoOH9Lf9mR
gr19NN5KvO21PQUk80jEP2DZ8Qm+t9TtHEX2YXrLuSER5pStS0T0Cdp5s48lvDu/JzQ31GtZaMNV
TneorwZI/aEiemkBHH6QYo2EN5Hj/TF6mHIPAcm18Sr/9jG+TTRBnKqQrl8gFTKfwyIq7xtVBWeE
hqS+U6+Wk9sqcAb0h57/Bh7EeUZg+pUt0pqEVMsJlgLRN3drj8tyVLRGCcn9GQzRsDa5s+F0gtvC
YZhHJ8VtZPG6vGtjhhYXjT5+h5rSkg8RldGa2PBHsixYfKX7gTLZOcs58HhA9FRSVTxnsZuM8Vkh
qzOHVCZdFC3M/48afIfQ5JuVtQKkqGynklsY6npDZIZqP/yeYjeRam/AOr8wVPewf0FvnImPsxWT
JISxQ/GdEuRrhIGtZXS1T08XM7u7hLoJ5vnG4R+ly3Pn4RJ+ir9NjNdbLoq4L9UlXR6dfGd98AL4
ICHjz2FoDJ/uQ/kIQILL3aUYgRDGAuZPaJuLow8u1kc7Qm+udPJIXonYqKx0X+2ZmD51ZMY6OprD
GgyqiStreTPOMnRAHyhD/tfpja8H6BQcllBdUBd+o8WX2VJNzPIrztoz/aJgxGl2GZhO7cE7XtwJ
Z+obkItu9qt8fvEhksNl00gy94DtyFDrwCDYj7CCW7iIA95Tezvv8P/ebGhvgXv1tPEz5wH3VSWa
Ndw5e3DusOLavUYn23LVdESOYHdqDfup7fzHM3WDwaeby8OrcjlcfSY8D4JkxafKL9wjg2fmYX5V
Nfr0nMCPCfhJw2bDHp7TUdvc5duRm6B3aqd0Q0HWNVqL0il4pGJhvX9MHrRJmh7s1Al2sz/wSIQE
TWqyHAoD6INyxbBdfct+Hr/ZpMNGSEIqxqrIWTvSP5SxxNraSBA7nLObok64fV632cuaGT8ZUjuv
dLMLFAAMtmfbfF5h6nmFVM7gutnnWLSZOMvW78pRx9JwdcLFb2NEaaKVtyRzgnXE384WtI6cdkzV
SW5LerFJoTYuYWVDxLKXGISw7eweQuF2ISmCtLNzQdZr5IeXKTs67fCv/INX/xvOwuZ9Qw4Sf6Tj
rw2qKpH+QTWkBwnvf1dA/6JPjhbtXHvDFD66oyExT5noCvc2Dv7pidAGSHPVQ3+A/f26bg7o7/8d
HAHTr53ooxDg5Cq5daCSD3y1kJwkAg7Pt1rNDd9U0Vf6XjZNsozY6Yq74OSkN6qe57Qak8zJoB8C
md25OQJZPewORcGfswjvjSdFk/ouPABpgbO5kl7rcU63JDDILB5d10Z2QDG35L/nOPRFv49SXVv6
BFcPAqe8kdMIy2/UQnF7euu69Eoc4ZQktmbMMrXy9jLjz2dp8wXbyyZtiyVqyrwFOl0PtD1o1m/x
/b9r8PEeqXCmOaFA3lwswOp1fjseRgGpK+4TQ+zUCdKCBlupay5164vmD5C1s01xXjxkRiAG3s7+
+cqbG5hvWqUH5A0XrYeY7imKJn/A9a0XvV2kWj3sClyN9kWVcOJyxH/nTnCPVjP3cl2WHwn2QQsb
c+KEPkcugsHX70SP72iEqJbbP5Sr7Au0n0cJfU7rYwoHUz2A3X+wghkPtpAlacMAVxofCja6JMmS
gpqHcD0zlSxcfXjSyN0LyfbklXfwpppYpPdPBffRdMVvwNkDwVL3ZFc6eBd3Zc5MjCeFphZccwyH
c1csjFi6rlH9Fp6Vqp310m4K6y2tibeh59+QYg5Dnbvwj0zEuO8UhNPVUeQzb9378ouMB03fPEJv
24V7crrUSKM5twURCctqb8JCQk5mu6l5VzztxtWqAP47iv2LDcpnhufzkvuiBr5qbNwJbx99f+JF
jhFmJYajPwd71LxIuKrC9r23rF6g1r5japXMspiW65cb9NOAtOxwR4qhIGE5b/M7vncwCxSYb65o
oX+98GowrqzOUCoDHSuKMY+us42xfqMIxPKCKGoAe9tDk8lpOZLdCrEVzXkIF1dcHBc5TqH75yxI
IwNPmr5Wi1c+3DTmjelycsj89yWPbmc6Xc1tRMJWXhW9DzEgyIWWWhT1SK8/pifX+DgDplrWvJ8I
VX7b/d66mgEU62FFIRRxB3whksI1o2pAxooh3hztKE/h6miqwfce8bnhnUZcy3KHHZyDgOjNcSsb
Y+yfsDEyHto6sIJxzelbrf5bCA+4F0XRvjYMm8ogoibabum/7COhxs1dTUS6K6lDl8pN8AKC21uT
9HRud2z7C8VXUrExK3zUmhlGOczYXNMNTYWHhtn9NswKtfS7B9ycYK8HbrvkU260z7AevYG+2d8+
SHdhoLJnrinM/CKogdbWam6jw/Qv8rmerIH7n4ZMupSy1TVAeNg+w7r37kIlKHqMbIgfvjbEADWf
Ipwohq/YKiIenzLo/22lasd85F9mtB8RXjMx0plSoU9b9EqaG2olZgQYKA+ovqyMwAbu4Ov5gsaK
ehyZIR7FGXex/ZfTmd/fK0xByT6RJGj3sOhWRPKo6MQddndHnQJn9f+EbSkQMOlbFvirFwmejH/6
L/2cvBrFSp0DJl5fqV9FHdygIsflIJRMsL32yrWFzZ2mNZu4lVA6VIY6NIL/iV84bKzRJXJS/Oqz
IW7q+82czmZYv9WNoldC+pod9ksKGu/8T+UPXBRX4C74H9yNXUzgvDy37NVJG7dyirhQHFlEQp8k
m+SR0mfXlgcO7L/XqMamb5W5XbLcDLCS++AF/nsSTYms4ix2/xfOzi9+ASPEXM9kPauEVdl2ysTL
PuE9Gb1IlfgkXhqlsd9PAdObaXQk+vFBRqcVTiWxgTZKShT+B1DsHdlQDcCBr/vc6XN0WkjwGnG/
AyCZMaQyvSJ0P8mmTTTQ6gZI/JxKr+gTukDJapj2Ka1zRqbIuuovSAtEoeu0JgjQQEy1gU5ISMhz
aovUWrR8gQFK3YCFraLoKjrByXZYi4M/crKDENrBykCFb494IAH71JoUrbEzFwbCkJktsyP2shbd
WTmaDon6v6C+Gl+dS/RYJ+ifF8LC70e7HbNc79Hcm2L5AOie2+EehwapqLcrIvjsBFoqdCz+m28b
9aiZt91e90H1kvVRmxx8FcgG5Hn5z4hf6Gu4KlS3L3hThb1ARR5iIcst2uURfiDEKCtNBTcy8Tko
XCm1cU8PceRiOXw1UtYfHJFcUqJ2q7PXeokqA/u1ktRu14cL0NQ7yspKGziANDV/Rscq+2BxQ7uj
kOZaNpCHRYORYj7KPVzh4t4zk0AfXlsQ10mnrgJyHce+K6tqi67MhJZJIB4IpcccPHsWowUn9pjS
mlXwBB+Dv1fk0fomVpyZ3k/HnjIoQ5PAAjWm1SBoWU47SN8q8W4R8qhQnQAH0QfGluexPDG33l2T
hn6kaz/4uILTPjT52g2CIN/YKzdlXsTiYCyvB2YO58YoXaH0LWj9BtwvBwLiryvLBMPFXbNSU1L8
qXlnU8jjNzWeCn31tQZlNx1/bM5iA+6LQCiEeVGOIs+J5UTWfFgm6neAJwOSZKtpidBLJCK+tNi0
sqY51Opkdo0/g1dh2wrme7M3iimlST7vR4JQV0emx/mVrlZFbGOdJnJcY2BCJSHC0nwJWId9fYHt
mfEAPznLaglEaOUVTAQdHY3VpGcgms0nvBeD8dHKWcH6qrHIES+eQzTzvXuSFHuSTB9b2nLC1Ha/
4DV88bmXbqZYhHlioqOF0bTxKFY7InVnd4yTlMR1F62KyVovd7vWX9HOLbNWn8HsrPqy8LRbXjxq
dwdMK4ldmUjmbrkQBwe3CRTREzFk8i0k68dvmYgqba5Ik19PewdekyS1IxjA7/uS5G2MkUguV2wN
mkupEz4J0V6pEBbgOcG1O3SkPwF5UN+CvZLHik3RgsB7L3daeerfXED2U/mhhSapyNnyeJJaiAro
abXRcmlKEJNFkXB022P2/TBujwGcuW+3WQtfTUxAjpN6zzjz9e5yz+GQdZ46R1DInmKGkH20pRhx
uRREN/+paU55eRyfWSlA/kiWevY6LVNa5zBuftyxlFiExUHiWV5GWCCFgwOOIXJ79dN3R4ynXQyM
lbU3EJqdcw+Pv0kUQe8Li/QWIr/r9OfpKyhR7clRoJXxmwIlp583KGMQGcfpLUOAj9C2OxXJdsLx
tA+G9/bb8ZuyA3t9auFNwf2cPRZB7FbooJQvme5gWSXRHKvkwOoaA5cSmpNNZWHG7LaJz96HZDon
KQpZlaYq47eax9daJBliVNbrMs3pi6V3QBHGq7VAiDH9fvwSbq0Nc3v8QGFUsl4UDerKrlize865
vE8a/Ub15Soh3b6mx0UilXOKouhtsvL8+M1LP3EUoptx/bJsosCMUoK2AAgRIBuQbHJCPCgBGExI
+ylR4GKkUBPj8IlDb0Yvgu0/sdVMzgytbG0k/JeyMb4K9eCxGWC26QejSeF4k4Rj3GqmW6NGlBZy
v8vu/GijcXaF98fHJfQuxexyJ0J6vcw22exX2AnG9X6GAekXuvJyQYwcnG+u7vUiGBdRjFRRFhc/
8d/9sBI9eqAA8a/nbt0aeccTdssW5+H4Z6WYThWFDqMiuAGSnDg88WiAyBh1HRY1p2Pz+bc2nJ2W
47LXc9WSOpJBNRpL3oSySy0Qn18k/PPzUPavd4he2YruAqEomfdWkFVYUwx8UCwo+vLdDD71Xv6h
u5em4SNdItnRu45F5285QEYErGCwf0IALsM7SlqfrOYsn/uhoSE8WXcJs26FCyxYzxJJwGDi3aqn
2OcdVmN8Xwpy1gEgzlF/JbElSpoD3TEm+A9kfjYF2Ii6XARxQSvZzCBEkoJE7pWYsa+2sm0uRLpo
Nd3YMk42Fls27GziS04Dox7yj+ADB0dF4nQsyco6T23R75VtOnpPyXJVPKL+gYhuMlnVN/bKVVuB
35Pihhe6bJwiETPk7GiduyznH9Sykobdqtj44KRFiCuKG7UYwIc1wZB6FhMTWczlBcutY5atnmFb
bkta/7KTlb+Gxbf2AWhi7MMgchZ6VErPAhY0geZPz+J4VfY2XXepB3L7e+gqBcsgSND68zHbwVSr
u7huz23IRm/RvpX0ROxtxrm9UXgCGvdjwCg/xBjejzDLZua+8XXWOANKw02axMg0mQpoBQ4MOuLN
7EIip6YHKA/khbVtkUs2PB7LkBAp/mAtkQnilo5MVQbp+TyQ8U3i9SFYGd9I34EtReO1MwsyLzbO
cG3I3nXBgdCZ27RU9jPvLD3FpSTPMHU/JvKgFy/Pc9r2fvQl614jNtzPDzRFLu29GaVxutmh777p
5I1Jda9nc3toO0KUriKvvYiLnjdMHE2kyc9/144CAQqZMdubgjKEdsBxzVExYDYeXce++tmlUoMn
8/0x6jLPO4+kLDFRKHkG+cVGkH8BE68l6JbjcUrrPHxfZ5d5/8acbSHZNdATIYnrP75F1vbRzaWY
r1zPD6QkVTHc2EMyusOkNIw3KC314X5LAqInC7mBxxCCXO4ROxuWz87JImmYGI4Drzvyap4bPEyd
Vt689GtB2R7pTIzFRC1D+Rkrqy2ShGqoclvqi0ItEZ4cmkX6MiC0FEndjlQ3IfVL94Sz1E8UeAZr
GNG4djVb6GCHdjjIjXDOR9jXtgTdRG8iLBcchdMe7VBaXKSX1fsXeD1DLp1VLuW3kP3PGSNAPKhm
bx4yWfoATwvVTBwumc2tHSSDj3hEs7pmd5PS7C3ddVm6MwNmuPj6LJXQ8zv8isqCAUZnOr46CJze
NQ88EF9dl0KAUlFPALKZ/Lv8Mj5hHtI2RRP4VC83SNz/X5+cKvamPhknD74YC4dxxhzo8qYgtexG
bj796FFii1yUvkFazbOTs0LW/ByOo76uCbI0VEjukWJT2zg1PzsE6srtTjq3PgwVB53GIzTbaLA7
XIa+3zVEIWG/rQtq6oTCQptVWJiPwqOkf7UzMF8wcV983FexKkuDSP/QZ8k0ta+u5oLkgP54gKv1
Jjqmi/C6ZqC7OCcRQHcptIr5YpCWraH8GcyahAr/Gtb8T4C+7PuoritcB09d89ex/d7yge8F4lFy
lWNWUzG5naRloV7bG63WL+ZEKSFmT6X+B3ltrU+gdV5BPr13w8i6kQzZ4Cb5BSBRZaPgCinkFhP2
sYRVGDNpZV6fbkbbRECaWfiu3XnDoO0nokDzdvENqZ3SvlFWmNm1JWbFRUezSrbSaR4qMXv5ozAe
6R5/kpJXfZQq4sLLMdiFGdLC5wMnaYh0lnE2E0MI0xOgK2lyFG3Vk50jK1XOHyeXfBhxHhP/UXMN
B4Yk89ZnkPAHHUDCSEpFNRpl4tnZChv9mhL4BZ6287WA5yoWRxDitjQBT/fbQq+gtYHU9qsMwsUN
LWtqxdVt5O55DuJC9JFBX/mffua2c6Vo2VHIcSWCYANINkCYrceYjMUIpW39fJyW/BCkCuqCGXN2
A3x7G0FCTYPeIwPAkLTrId2MQq3DRJmbrBLwR//dbe7qOufz83AnIA9mc+ispWdOZAuessFXG3/U
ZaQEwR17iTnXKikAd/HbmpU+3qLmJI+KLjsSz1mxp+kGzRMip4MGvulDTOCONZZlnBtmFZUS1/FR
wBNurz4IMyLFtLrrwx6DTbJfI2n6kJVU2RJMtjbXWGYDEnKB3B0n84cpkkauoJbZdvQBldr8G0Jq
eY7Z6UtzWAEu1P9y2MI0nS1cq1KvgV++wp4k1DFVMhAeUtgyLihY2RW4FYrPGX0JM8Eis1PSFlEj
GUDcWovYZ0EDlJvRGvAh1DK/ALXVyK6/5E9Jha/jYXBbtNJd2aSHi2+JgLwOXUsiBRujUyQLWDqL
g8/b9k/jVJCB1T5fTeHhg+nPpyT5KM7YXFixnz3ToQmS2lQcaGijQ4e83eWRBG9FDSBVaj1EiJh5
cdpBeEe36qF7HBB8P51wzDX1FLaYORZVNnQiI4TgGUk0klPJasElxW8HhRHVdc/kSsCSqGNvtEFE
uFJKBk9kLarjovxO1CphPKd5W5VbRWyrkAi8zzm5ofi06RLEag8+pEAZtmKPtc3IFVxlSNuO3/AY
46RdREKBKnFgDKWBw3KLdv1CsRWP5Ai8ODHe4TWSN8mU9+19m4I6FlxRb1jENk7HbuDeC7ImvyKT
S0h6bft0H60+XrH1LSLRkZxSj6RcRCHUUGyNKzLOampZIw+0+AVcTRe+slv3DxX9eUzQaNGWO7Xb
OjpE7xkB8CyohxeZIh9DOg3g+L5YO+x+uijtgZqDDRwxPBIIwlAZYbkvWiYBAeR/QaZH/9zRWEuJ
QyOXYPCQbQLmncvy7tC+dGEagqFs6Bj+tUo7ELsPBjag5Xj8EcVqyjOJwraWy1tm1KJ38/CkBuHI
cVsGtBR0Vxv9PTP8jLPVomQj6m0zyQVCBxMIgJg09E8zPa4roOf0oZ67hLYNjCL88sojxAX69hi/
Nkgob1wJgfHUCz2vGR88UUftt40cITedHcF+Rof7lwAZ0ucMCmkdQa865PC9SzAFPYcEOUA63mkJ
F/i8+6PCsU+bFttrPvcp/hX1ylMzltAYPA2gCUdtvh37dCAFpCiY/S1xwDJeAmvVALEgyNdnLVRA
ZlnZRhIXxylLmRGkgrdpC1Rw13lmfvB34jvsSx3V0eUrYSPO7JjKF8DQWNLf/ynj34QntOUJyrSs
ho4TemKIIihDc9/hpajixcemupiLhRmnDF8wxjOvhYHzkumuwFgdUAEQHH+PmxWMdBGnUf6JSIed
oMxHGmqsTlQeA3lvoKNo1Kd1SkB4kqLXeFrRHH4my1TR1RuTmBapM7jFIw2rHXHruix9mUaZPjJp
y/Xfj4zCPcYlYFOrtAJeQ48kO0i4WTIe5jGMQPNIVR9f+zMR4tPHc3Q97HQ089yPCyffEMijyhD4
By8GDmz7mT6hPKLl3Nxl1mUK5FrVPRm4bkAbk6OoIbHduKesLjqvnhFCj+RWhmF9ZURM8Wepb1GW
TGfIXQqCIhKOUudIaRm8+zRgja18plQmqhG4zcrQM6P3tD4HXPZ741HaGHNbAC6dWFPt9IP/TW1x
gCiWWzkX45caju0+2h09OWEsg/64CtL+8OTsKtFF5Jh2AME0kuU7a0tVdtraGU1zQKmh8MDLSs/o
bOEeuZ1wZaa/5grLDy/5xFnupiGXlxdSPfq0gZMqT4LywpooZN2sYFwyV15PV/LMYwNIy7151qon
rk+VI89v0IbdrlTqijDC74qW9JgYaHV4dP4zekA3ALH5HYTQr/ZwajFr/KSuTW87LhWfAMndwGry
NI92gy8rTJkXIKlyzK32T6Nz3mfx7Q14OvHaIEnlI2WkCd/87ZGR/li6kbod3xueZk/8NFK4coOd
y4LCE07XFc3PIr0p981mfsCAuz8RR7aZYfga9Ue04/R6r3r3FxqJNMPd51W3B8mqdmalsXyXB70n
wUgezCUo1tGLNUELtFybZt7jE+f0Xam2VuJqbq4y1v0Pyh+/l6EnUTyXlNtmqWI1eN2QM+ysTc+E
ld5H8Vxf/eiN5sh6o0jg8vLSBeBeCkDooKYNBXbMHWYSIYMg8op+yK4/DfokiIG3We4A6KG8Xr0n
WFReuyxKiNP4A6eAKQRgmqcERYUb4T7i4P3rDyrnEyZ4sMez9CnKXrjHbPIZ5Lteb/9d74SyP655
4Aa5eboRSbrJ0LbkI1UneqnLR0phRTtqdufJvsf5cfVLx8AQ3lNYgzkGMMUUlDV+UowE3ECvM0Pp
LS2Rla33Q8P4UAvhf7lLVTD9PDyfIrCnbpnlt70G2/ACJN64c5UaIDqVjrJ74FfsZYd8f/wxQCYE
0OPrYyvg5eVqAuA5c3UXvz2alEefpCDU1P5B2FbpcANbesD6xon+IFvaP8i6NnFFq9EVbuhMuQNL
0CpQhW/RYB6Yo5GpwJysIeTzhIhp3l5jew3TrYKCYpvmsNBKfAqofVXpQASBYxRLwTmTC5ZuWuTY
/Ay7gx/MODoTJO+l+yjkojpUeq5zlOsMjLXSOJAFu2lhdteXisWiSH6Q9nEOC1ao6Vl7dpHWjYU4
i7SVPAeTZ5GfYPIZQuAaa7Md7cKUQ8VwGkAJQyvqlQz9tYHp2707Wq29gfWo4ipuVnq66NTV2QUb
7vXzt7V6bLvtmFKFy2QOX30bYeQciHPzvSyHn0LSuwQ28iJNSNCI+V1/raXz791RIStuLvS0q0mE
cFmhu5i4yIJtjov40SAVHwkzUKp5LavUUXMjyr5V/Ts+20RJO8Nuv1KPgQ3PABjdROPrRkddKKR6
dX9PTbgSFFLlFLgVrJCtf3JsJusH/ohLI8c6aIFyt5HSZ20wjAp2X+6Fn8GbDHhxhpygLQNQcS0o
Jk6hwokwonMztII3SToLj++NbGQxMaseRyE/GiWXFd+mIh6BDeQd6zIau9qKgcKxl9IAL3n9HlH7
7cKgk76ULstABF2C6jw+F3gvm9DQO7ZajolWiIrzFI/+8UoYmogf+X5SXqsyZf31L5tooWSxK6kA
hZHEijb0+INcPIyiYWt4ZWH3pR66EGjVOABMqMB6D88FIm85Px9aMmnA26bwp3VhGE7AoEXDlPwk
u4WBanQoFQN8rB7aNJAuCfMTuX5bkODcbV1va9lpk2oyr/VJyrs2huYjjrJJaL+o3Ro7shpIZ4Q/
a22UDbNBg/abTSwu9CMaEmTM075uGbwk8fHV1U8zEZAcaInepuKDiOCqbbVcSyUhu7OCB38inzaN
creGP5Qr/pprnDkMcqTr88r6vktE0XV9xWCjOfzkv0DdVD+dZ9N8lm7kOmQDp2sIFwwfxPnecTNm
S4M8BR4pkjayl+Jz1KI4rXqZtl8mzQAbK0E+BUpiIThoD9n9UFw1T683+PkfTRyMXF+lell6n6J9
B8BSudcV1HU7zHgHJATNkmrrbRl09ntU3jcMJPBMMViVcPAombkpy6DFkyzc7MUifmhmzPVGO2hz
HYLf9h1qgqeWOmjAC1IszGYnNWUUbx500Ys5MMJ7j3JXtEoSgbYivqtxeCRaUopU6ZJiIkTxfc1r
zRRGznxj5thpLgA8cMYrTt/KRWJeRD5KnmGIH3a4JGPoH0M2SSHlnc9Qdh5pkHL8Vgccy7pGEKJ6
WvtrgHYiyiJaMtc34q/XTOk6dV2oEKw/xdRveRNLAKWb6Ygy2xARZHmCtgnHBhPvoa6eDhpRfetd
xYdORPC6xzsj1U1GyGeHohc0v7kDdVNOBd0zOC5ZcenZDbz+TfXO3GqALHkTxmDiTNldRZzk4bXB
Z5lMwhEO2oRw9yFxlf0cwSgR3ngbyWMNd1CAs3GRjon2d1F8Pw/LDCkdTOliUyWYt3ofvI6CSZui
MyDlSm4wB2GtoyYuRN4C71kpsaol0dOdfyF9XiDaV4F+ryCLj/h0+r6pZppcnDAeIMvd+42OQPlu
VMCiLukICwwMJBX4QhFf+bwS8vTzxN2UaWQiQ2pk3cwA1NH+21CzEBbWV4OvL5Lj4njKge5duliq
/c6Kb1Gwd7ksEzh2fSlJvBHA6V2efaDxbSEtctd5KHQd5+DQI1/bYxB1+Imfh40uWBoftQAQ5JZO
JnFh0nRyUcTF94JPnJBvMAU6cDkjp/y2w7lpmMdShjvaGdqmbO1Ka2tE1vYEpioKRJL27D0kGUSw
8aLXTyBM++b/FVz0wkFU8VXaIXcwEsroG4ZdOgnOaLxHlNe1F8cLC0rp/+FiZ19BXzUXCi/8eh7D
k11U3KEukldhLwZuasb59AGMnOtQSK43X0q6XwtNmSTxpLJLGKMU10fsKvNmmQNTYM1EVlRN/Oh6
volVYk8fZ3TIO4HEHKcnNoG+PyOxfqQzowSCCCP1qA7Ch6KhQFFgCSoFzi+sjqgYr9PvMg3twHkF
lWg5E2eTXp7e2M5fDbl+YG+GOU5tTwIgvDrUX4zJKHdft2/llPNdRHkhg1Bo99ITjLlw1I5XWslu
aTZxzPOE4UsOFExy1K6TgLVcxCCdZaz7u3R8NOVfvS8TE2UveehT21EU5LAgHYkwTrZmzlE8LA+d
rTW+EO4KiOSu9ixBW9BQgy6Tttr1sy6yEf6ov51sI0QCWNfrgdhZ5dvoA6Od5+H4z+jEgnC9kQjb
4Q+6P6kdzpS7KWF29HngJuzODOuSrlyNCgZX9ITwdD4DEM7LW1P6hy8le2loOt3ZylgBS7N9Y2o4
EfvpjYYBAPzbLvCeRqRryscH9OZOT8DKCMWrCpz6nLDni70imbNEPIbgfohsdwoeDjVClanY9ggW
YnyPWxuN2SOvWlRZW7w7qb0rkjn0yf8iwDXgKh+Zgddnh2TKPKq/so8Rj16mHY+GnKkFqPCwqvOI
i97B4ooqgrpTpJEX6CLDWJqoWIJxZ2LhiaUjVXP9XIO9/0Yc6CmfTcufMQ4rIzjsJ5paFAkOHur9
U8efVL0lKOT8rAVSRHMmHwfFfIItoARWmQjRq4cMrZFCTeFk2uhIjf2DS0wrUf2WqMqJ9E9HfVBv
ioNVODgvXK+aBcppf66tUpcHycp2d6Voj+icYBhSWB9XaH20qh36yiwO26r7ocwjXpREzwFY+q6S
3cLZWQrbr47ebo8K3J19j3xuwVFr8DiTcYMt/1MsX0JXRZFjJIjl6SDrKcodmgoO5yp+eA+JiCJZ
nLZdKkB+Qb4RJl+yv+8VBPjQTT9UeBJ0p4yPc5M908qO+PgDaWjiH6IZ9eLG+MOmIUAKJilwkVZu
ZYjoAkccIR+Q8Wk0KFL6U3SLq3HSdJQeqSkJ3dSda1iN6yAjbOh9CHl0WBuNJDRy1pis7M60Jg1D
CnBzbg+OM/vgBdD1Pj7Q6D2bHz+xyHNDBvwSWvkng+7ISq2enLjHRM70lYxh6wuudyyehCn8S21x
EPkud5I51ImptK/S+4cAFVtmgbX/CZh1RYvXE7Ut+XP5JBiyuarXVOd6JtsVvxNoFcqyzClsCxgb
BfQQpoJ9a+dSyEzAbtmYcE2ksjAg3bVg3HKXeotjWA0Yu/v9gbzrSOFnGzNpI53Z8DvlSxITY91U
L109mKZ8DitQC08SWlwZrM520BLTS0jMhSE2X8g9JVdPhjFFU3Si+Bdit74+OAJrc/h1lRxqeaXz
AVS+nioW6XjvtGwpfB7u2mgHxeQopHveQLzjv7jA0zlZIhb8qPu2/5oGTRjNLQ8OEMrKDnZxfZ48
68W7qI0e6LNqDogrVCsSnZwC9MTgn2QFsCSgCMn/kLsqLpU0aIpPTldRNmHc3cObxJPI2ZBGIeFk
ikRiPnrVnLZtSHuNTVuvSLH4up7v54pe7IhPbrXCgZl/RKPvcyESb22FQl9fz/TfnGgY/QldAPMB
Dq/uGtgvHUjnESt6V9pSfMA9eltYm4xgTTKKLAbzIqdhr1uFAWyYuM6KUCVEY8XO3Rb6+yTbaItZ
x+pUqYdpj2onJjzGcdciZ2gK/AGpgPsJsJfj5ZW8lfUcVlDIFzTpdXM8Ysgp+MAVxxIhYv2TKGZE
ZHYBZski1on0+dhD5tWO9vLjJ0zG2V61yvkhGfztwlbZ3wpdf8Ja8YJa/gw2qL1muwEs2z+/eov2
JyeT9DDC2B+maQftA/nIkUIHTXbt3OUBZakm4JUZ/6+BlZBAJaehTRIgegrzAu4wjzGwtzwbNBtk
VIPtUFLUx6VYkzLPVyGTgehDqnA1x0dTjXQnZt0bY3iaNnt54kZVztfzStpE0X72GO75mEvRT+tt
N/cyc8Pw/8LXaeo0n+961zUn+o7jYchYSFve8xrLF468FGHTeNp3aR/93tY5jU9QgN4W/1fmZqP8
PxiuPEE4bvGqpH/B5C3b++E+bpKLcHQB/YYGt54kUYtl3iHG6rTTzwzpVhMQRnIJmuoz/fjS0wax
VSYRbTCh41jf1F0R4TH78GVxFy2ZNl0mmmyv2AqXLY8yCloBlUhjIss9KEkXnOkCCi4hrd0JeNBC
MVDOKbpBS5d8NuEAnA6nn7kAr3HR8WqNfguF/nbkXKNBa2nDjAfX4KQPvJ7iVYykYa2OgxBoI6Y+
arIRzYcHx37ltxVyCsIy8ApxLKO3bbLJrGKT+GwlZNniX4VntzuJ3aPwZwQEj0+qm4G5oxSpJ5Yy
h41i/EJhMkJhOWYslayJPIhnlK4rsp2fT0wd9MKhoOrX1bmtTPDixbmRBZNa6gQcP8o3/buCAWji
gU/MbQ9YRPAracuTFmRdGRxbf8jDhsbS/Ehj+CJFJ4xsmTgtFWDanfWw2wKaYkIwmQEmN8v80ny3
sMJ4LxDdG5N8aF8iEKim13RPFY/uz6ajVNsbmJbG5ssOeDx7AcFO8lkg4LnIXbg2j2vmGP5S1AWI
IE38bJ8qGU5b0LV/lkrqbKQWLKfLcw/MfeJ1AMMlVdREUerCk9QWyYeleGNFNoMYxi4N+jw+VcXv
TlVdWNWOo2PAPsaXZugZdoT5WAnhj3ZGho73b85twJKS/7mzHyp3eDQt49pZMfnpTWTnLyxb/qO5
OJjxvGQTNAu/tQbi9BKYKG4GC0DT7FY/ZijF9gN1iJtcgIoM2kuh0UxoKO9dHxT+8mRNMSAkRGjT
sfZFdLusU6z6pRKYSiHhenxhA8HX7CUwoeGz4IWvoNOT7OwP9In31MwVatXgZNCzK7nU2lwjCNrW
rmGsCS1xrapEQmDczKVMhYkjT4XH+RrI5Ch6iAH7JByJjclmGSCkyug7jDZd8s9vDwmS3dE4/L56
BwmghJ0FRsNuagB4xG3Zi2J8PlqTh3P/v++nIlL1TFa8AOTi73peU0jgIvh5wo5Ygba20RpqS3pN
lj+koeLSNXZz739KrGilC7qvkZP3e0roYVIWU95MZ8dcWNU7KT3ZUU0s0KP01rq69RgCc1B5/EcK
S31Gsjt41vh1LITQ+JranWOOyLWjimKtB6x7//9rc+8AP8FZdNt1Ybe22S+lCPnKKgYIr0wUOErP
NuPjyeYLh/S0DfuZmTM3Pbcyb1SHE45BbZ8yHQllzG0nmF03utkAuXCFq4Gv/VnDJHozpHc9krA0
M6Va/dpyMrhGfKSWHDX+Mckq+q64pdVuXUXR2db+dWe+Ck8wNIOVxwCtBCYStD7ovZx06bpMigFC
VPI2sqCzXDZKJjr2/3VDgGGYOHQdfnYcxh3tXzPXQJK5mEZfMrK9WPy2YgTn10ofG+iTWlMfC/o0
e2WCHMwfOL51YaEhSyiJOWarR1T+AV06PxERtyk+LbUheDm8ZsB62lyAJ3NUiobYEqhwzNXHYMLz
HKGTg7dFutPDqj97KAPc8WE5tWv7I3iA46XgR34rhkKxy/lx+ElNYPhH75NQUpW5/o2rGQo3rAtx
5VGRnPna+SDfZ/0BtrUrHfqqGSgsie2BYEjc/P21DyUqCxy5CY6IOw4xmVFemCwnVv3TjCvX9Z7P
Vsk9ZllJO6aYUOmgX7dQnspYIJoIaa2nrmN18j39JcBuc229BgSd7figFD1Pgs1r5Xed67aDx3Tx
uI/Tk9TZc9szZXalUY0NIFl20ZfIOwQpBfLsrWgQeESBJ+Jgs5wol5sju4vDJu5K4w3e26Lc5lJy
ee8+wnOWBBW03JXZEIV/L+nbl3pGSjOEleWq0PvC5IfInHcGWT/xXZsFhFYe2IOD4W6B/lD4QSVb
/4GjHeB7Lyy9rjqOp5stNj1/9LyqZUW3a+74UYgcQbWfe+ysq9Lx57D5TmCa5YCYd//TmxlYyG+r
9OEftIv8vOdB8IDwjmAaW8ct6cimtSSNcbJIclrkrd3tnVXhHGyvknHaGIX2/VayJ7kth98yQDgg
gqolKx8y6qQKv3KHZhqkSv3XEWJFdWDpPwnE+ogIknJvwldklKemk19M2UO4+WrM4ulYMT8dmj4z
7oBb5snkDnW+jX3ryTIBvFRw5rssKru6jWqOIiioYzhpxIs8zQ5TjrjqZz5Upv/M+9+XsbhyncoD
Xub2jF4J6jwX9ZaJ1c5RJ8TvLnuuRpV2iYo0y4vkhHnJWGfb+AZir5Zm8g7L3mvt157yn7dCfJY8
RNMAugQVHx7NBFP2uP+gH6zLnOL3o8jk57wGgwGMrdmH3PPeuZRbSRIqbndBTk7Uv+1aQr6xCUza
wutEbXy6/lRDQlHAd5M1rdTJNZGV2aW0ltcAjPe63uG1Zb/DZ2yLMSLD/ZjMkK8pcWEKOxUT8qXo
bplIPSBVfKKo8wWZEprI/1Xls+yCIAN2Y994GxJWX5ebuog2Yfa05C+JPLNV3RoEhar+sN9kfNb0
ht+rhMygSsq0HlcFuz6ru3QkSE5BtTbY7f1fd3EHoGDLQPgm/VOTLYzaDR7ULR504clRznfsKVlJ
S8H1dK3rKgAMgh5cc0TPVotBtrsq3ouTTfbxe0f6ShNdL70Kz6v+2C6KoUO07qMwcG/cnQJr1Hir
bFyC7h71qsshaf0806fA23fL7WvFzh0aOzAT70hutHTuRpBwmRToSPhxOQmTMYlXlBp5i/Q42m68
jJd9APinLaRlAwuNvGmUW9t4QUZn6zfqC183fuQS29vTr1CPcOaVCzkdQayj5fr0poE5JaO4esXC
H6TrTwr7FLrXVlLDr4y0nXlYez8uNR8QPOEuGSyPHD8WnqdRpMSJbyT7XCfNA4GRRKDH3LkXgC53
AOAgbuijxTTxUnpI3DI/m5ng+3IHocgbv4vLClKBnMUj8RMfvZmBxiw0BeNQyOlKXHHT0/LxPaJT
BiI3WJSv9d5RIdmBQdveCgalf15DapnfE7ee6c09BDO4bVp7mrwJw0rbkgWGuxvB+sJ85yU0v18H
QxrGr9zZIlrVqr1UYISUAD9C+9oZGskinuKSYnj3jEoo+1lD+X0WTHXK7DEpSR3/RHv4L5KX2jlD
AP7GyI/MS7DjA6ehQGYfQzyMI+NXl79S8x03IRIz+6yKrUbZ2M/E6mBsqLyZz3W0xT+R9rxPHqUD
qHFW+P6fhaBMjTZKxb03VHLUw1lkPHteFAHCQHvvGt497lxZEcW7EMiMDNkRyVTJs9XJ19DdfMIh
1MCmF9kDgPfjkNBHfEpwRsF37vumVVUixIrqHAlxYh7uGulFl8PP7fcx19keqzgmxTLE6Q80CVb4
CGq5YFON1/uCN7vFJ6r+G7mQFBWb0Tc8ze+tvQPzWYBCS8vLnswr0kvbm7Q+A3LHD90gYuzXG6QR
2mBcTzTG966H77w+0hzshrwO+1fOCOWlL5VtDlzPVuBIfKgb4kJ6jTGRRaxaxC9BT36CRqY/ZABZ
WO+by7BXE5UY5fhC51xWnGvO+0ZtMvFQ4rNZpMvozIWDGMqvMzflr9vPh7BWmDuTGeav/mbc4QpH
NR0zBlPULen9l9TvmLrN8a9GU9mRT45VOl7wmGfYJxQOgCaaVTUrXh9Vgc5sQYYy1kNzi7rBk+ag
bMGLB7IkXHxzVlwN8Y1tf5x8OgGtoqLPAlh3D/AuSU8pLRyOeK7lEUR7Ue7v6JqdUPGs9VLM268L
HA54ywh3KTeLFaIXqE6bA3b8KIFT5O5sW83Frp63s82df4lA4rerU/2VsIDkATX6uFn4mjCabRGz
uNaenLWm3buMvpg8M+UTkevLiI8khupzSayrmCyaf9ETabmZxzcmTU6gz3fvSZUNY+SZI4tOPGHX
jfgHVoLXk9ZhU5gxv2RsTP2QRO9bieOe0wk5Ofg7Z3R8GJbaLeiwoFul06vIGpOHnTEF7KozMN8Q
BpTT76ELdkhClV2ktzuoBP3mKqCC/NmzjShA1AyBWNy3FldtGHyzFKuJwtVsd/hMCuLNHAuJkXgq
n401U/1ilGGNyICwSkU24VqNAdGNyqUw40aLRvfunvaUH/1ZnhiOMXDjjgxmQ520Xyx73YMxb6a2
ucMfVFWZHfc841CaTZX+xQEW7UlH3Vx+X/aPibk750yGAkie1XnhwCQgHmazusOwKClz8elH9KTk
ehY0kEP5cbSkpV/88LgJ3NFt//utr3xRvfaO7yJ95/3vVpLf0vjd7W12GYHGHiH2t/Ex5zfvdzDL
5SuYqGxegHBzZjVJVm5HiSHrS1eMrpLnszSbmyWwAJobvV4MvFKbaqyA10GLKqpAK+eBGuSRvTLx
xj2I9LmCmocHfZf8Wqp/wwkn2W/HxNPF12nAvFyhoDPz8Lku0l6t0ymmgmCvqz1BYAmpxydDX0c5
mJj/usY5wphH6CT2g0jB63rLoqZHcpMVCnfARf+ylp3eDeBNg4499mVw+klLfDogNsKzd53krF2P
db4Xd9i3acrmEogmUH3zPu25CZ/17fAcTk8l72JPZPBU9G0QRVAyp+xei7xnmRf8hcr9U/Haz3RR
ZHVD1bZlBW1ow9T7WgMVqsQwkZroLOyIEeOPayw2WD6Jkw2QB2Yik79/VD8beTE5hG9aR/NaCOsG
EVilzruAeM25SDtzd+WJGfa/PHWpmfLIrIWuRRJvyn2rDyvQtjxXh+CnUCEOu9cUOFkBC9yecv1D
43IFYWcZJEnXK5WpB6o6Rc2aEJarcLja0PdBoO36oY6j31bWjuYQtvFI97Gtf656ampH1X8cJbMW
X1vwWb4VOdkDdWClgmfvywaP8eAark3H+Qgbg/64lUmxJcJU0UYm7CAfkoD/Irrr4/EoQZlDFd9t
urdZaC464FN24JVsk7RA2Hw2+++ihNm3BhdhZlaOFbyuILs8p7EOT1qLnbisgXRiDz4eLI2jExnE
83E/59o4Y/7m02hFPY8saibO4xT+jFeVVAfcjB0D2NHQkfKTnHgoSwKxlJFYkd155AvCTbGEWJZs
sM0Pn4eZ0M0zyC4qWuh0cZh6Km6Z0l6f3/RB3826y81JXCboZR5nDrM7QXGLWQgypHeWHZelEgGV
528ymO2E2uk5bwytvM6ftvcpRE5BsODBsjk4G7sMfZI6B8F/lOb+pp8Ol5fpD62sZFKMTzJwM+RE
O5JCp/I4J5PDcE1XGP+gRfwSuth1cT+7gcvoxtoY5fPz2fOy2NSVCcjvEjRc1QVZ2PawPl90GwzW
aKh+GAePNKJmJ6SoeszmJDAqnH4uiHVbpxmoTY7UXw2O/+90YTaqumvmUM1DbsuPZ8+5e8DlwwOa
gJlEvXQ9rxV01DIXz1ce4fq6ma2kt1LO0W1+Oz7/DImOHOZD+siHzKE95XMtL6BZuc2yUp0As4+S
dTj+PjA4PpcdN+nFPs0IWMt1dqPWP3cXQMSm1jEuuYIn/q7W8qOPf7zjqxoO7Dc6J76QeSWE7CMv
WxyTPeOZvHcWCbnce1hiW9f4NG2HhMfMPkD8sj1ycvcmZg7fYTvL7dIX9l/Ya27+qzDlknu5ViM1
1YCl/SOJHwWeDB1WUK4QJ1LOwg9mF46Og5iFcH2xfo+/RXshLWjF0lACNvq6BWYRmb6cjBMBfluf
d9X8FRUS0Yj5O74ACGduIVG+ejBsnh80t3wBMjpqB2ono2URhVm5zSBFcheZzujSmRmuc3kj354B
j2G1y7KpXyS6y4tx8X+VVHCkyXDzC+7u2rPSaYUAsa3O2hMUBx65E8uELWp30akNOquMVaFGI2Vv
SaB4f51NM0mykV3SFsXPkseJFFqix3DK+/NWEjSfAOdzUk4oeLGLgTUzjv5tUxBSIqrU14bznPfY
O3u5WLB+0+m6+3kJH8/FNsnkncgvq/iq5QCLGiuPyaO7zsf5S/nu1/PaNF/YVuvHv9S+SwrT/Mw3
m0mowqYsaiHdGf+4hsa4HlUenrYzYqFnqHWz6hEK+YY5USQ8Zk/dgMA6WoFJLeSEOaFWRXjbjgqF
IcSPJZxVzeN49B1lLq7kg/L+4rllObgjaVXhoQHkLS/+UfgS21Yl6SaZa8d8CFy2R46KYVtIqjvl
yNVWw0grjEhLccb8Il+Bs5e+tt9TWWxNwJIvAifbsi6nEyUUDLeZ672b5JxDqBQr2beBWwYhxHEH
4JsSkZGn4gwRwlKX+O4pOi8rtRVVaAPitjUDzJO7VoRt5FwisHEE7ljTwuCcUg3gfcuW9wxtvQ3V
aDWfjQHniplpLUW7uByGedPyMBpFXTgZ1BZDkqegLk8nEJsvOT3CQ1wmac9vT0jA3T601NSOABst
wnw3Scn5hZc+Hb84Im2rHk3nrEsJVCqMj1vMs3fMy0MXSWIrCwxdhgHfba28nw7LFqfh9WWlqauF
9vkJkT+dRBp/JiGhM5qnMIji2EPzP2hjwPZF5qFTs/tOXZyGCZ8GiR8D9mF041N2RxC+jQLIAZf2
XaZl2PL7SVpogIIC2LeEu89wBl98klAlekq2s1Ckgv7pJ3eqXZ9b4lgBnp5bLbD7pk4h1vAkZXgN
UOVHN/ot4webQhwjYsPs/pNlt+wqZaopgs/mc27UsUQpu9HG6Pijgbzcyg0rsMdHvfkuBXQFy3SA
c41WGyhxAuKLU7WoKAgg/N/4hwI3UyyibH+j6InIF+MbWplV58PQlBudS22JJoc5FRo6TPN7ykX3
pp5HLXeezGCvZuurhzGA7k3wvAl7rGOF+U0GjNcC/fV1E6n44BGZ67sW2KZcuigklQzd0LtPn0Dg
PrCcoGsnCBuF6iwGltrkwK361cvspqjPJHdzTohcpacaVjskNDi9HoqAGitsD+bgXje571k0NR98
hmv5sIHXsmcONcD/Lc1ddo4uJy44oBmf/Af1H1D7O1BD2RoOonXs6dACxR3BEdsvUS6xmtyur9dj
AptyBh/lrp430y0I5GzwRO7RMAM0nMFWjCMvLDRR+aS4Ctv31skKzwyaeU3EuL++vnEFNxR6ixFK
EjCBrQkY3NHmr8gE9Cwbo2bwJAxhAN/G60ZQeglQ/lLXh+LDqfVKrNNrI5K8xa1cVGXwsPT1AB+Q
wu/xU8GbLxNHQA+waYmZeXKEx08IUn6fcAav452502WORejk370BuZLA0ImWmZRSwzzG5lQVEEkb
s3tD0OeNxgdxT7lqw2ks69I1UIZuglJTZibjKHGI4ggvwH4TBWudT+leeOxhCw85/RiXr9pT3Zps
ErCZtOxDKiSYBaG9eDvJlFSQcRNEsvOx8rNL0ak57TNYZ1of5x7xmNdjS6uqVCCL6PeY5nKhOtLY
0xe6QYPPk8RUXQs9tt+kcpoC/Hr2aihoFLeJrIsJ5hgwYPztca0mFOHcGBo6ESMtF0bzO9uWXfiy
8gkIkJPjOdn6DQcX4N79qAYMBR/FhqXDlCVRyFRV6paDpE72P/4DYlp5f0vSfJ7DZ27eWYpPmD9D
Jm4Wq3jyOgYl9weZPIUJpiBUyGmMSsYdb/J6tUku8ZwXFspypCOigwKg/TTEFfOu/TkHV2gLOrhJ
qdlVfnuQCSpQ0i/bw+dqAlKStvp2Nhnq5mijDVLi3NPYTMWi8Gpa1V8hN0tiI0nzEnA/QY6Vngmc
1WhNcBZs38OOGVQfB3xRwlDjqwXux18R2sMU+7Qtp7VlsUiOrWik8KQN3dXJYM3LrEXTDewJlOyt
UycPULwUh4i049QkSqapgtkS/wHEc7nShPgkEBlfBWyMUcCCncrIT1r/s0zEdC7uJyXMtxrntoy8
MvGWJ80Hs1SqdyfDi5QQdGSND5QfP5FT/vYvEn+783V6jVeJ1hl1id5egsrWLdbUSEBo7V5tG4uO
GIL/+rj7iZoq2kHhEFVBSmT86FPbGj6iZlTzTvFhVKZ+sOZTK1F2Fg5nY8b+zrws/yRQEueRyFF6
vP5jogBkHjSVPH2nq8kKAPMYC8NV86c/f/YoecA4HoXOtX4JuY0Q3HWbPO371wwpUd4tgNaH6k/s
TyLu3AwCnyfWICo0OPrdSIj9v746da7mteQMHMPzcBSymgfWPGMoNAquiEhODuhKZZwl0Xqtm9Us
XFo+6tWfVAdV3F3fR76oyoxV6YKL3RfW6YYuC6gcEq55Sb22rtioH5FoQ9SlmQmOih75/uKm+lDn
tEX9+UrlU9e1WKhhC+F/4gRC8pnO5Dx+OilCWdYFH3ttoRQVEo1q5nyZEN8tQC6Bdo6a4cT5V+AD
m4CD+xZi8wm07uzhA9nPhZbxpPvJYyoTqcgmCLklulYvHZpkRkkCcvsHv/tlK/ZrZQ5KeHhGjSxt
3sxwbfWM4ivQ5c9X0UZ8/IJYPPoHGaC4/1+r1L/xlle7AQqU8XTBAjFq170bw6XR11p8qZzkKZdK
L94KfEKgvYFlxgKMmzJSemKD6Y0TK4tZygT7862fkWQQecbuGB+NfRnMn5fPNFx1ZRoFOTKsMfK0
PJLKwIOZ8atKF1V9hpvfE9a+r4QX1c27R/koq0Rgphv3t4omJJbQN7cl82KdX3qc2P0AhMKZTqBX
wBsm68Ci6KB3pFYw9ObsvcPpWPPcNDQJDMnUXId4iaPE0ZlMn7l3rIUPIIBaaaMrrxr9FRCUmDIw
XbWp2DOxkxh85n6ElGDQXo2xPOgSrBE2LNF+rxVAmdhg6anG71auTBcWnkUM1lkRB7GJSugjdiPG
k/zvW2dNo6HL5SO7IWsAQdZxzOL5IqOTbSjE5CUSbHntCJL4F38dH3EMGZd+ARQt+mo6c332YTB1
Xm07oVYiFR7+1Chwjn7uQ/7XiGmwsRJYUa0oNPEh4Au50n7WjF6N24bs4aImYzL97j7fyLnUKhl5
ImdT1v1DBD7L2MIXT2lJd++pUvxOwAU3d11PXKAhcTmz+texNdoIdXlOsiWXWOCfbDlo/GlKqR5F
SkrkzTutTMGU+r5JsxEPYnRPblK97tCk5cdFjetknsqyVzKuWvHOvK3M+hWHk6WxvDuPS9wOmLH6
1LQTcS7DOgSbLxbNPiJ4WxnY+CUE9RLj0vDrKzAsbpLwByjCuzGCJG+NuvgE8IOHjcNBy6KelMJB
a/svT65Un2DAHeXjU0cN7Fdi6KbaMX0EdWfPV796nYaVjYx6wuyRISV3WU4KKrpC+R9vqlzc0HSs
4z5HRT8HTHfgs38RArmydw9D9czwiEbhw13Do/EYuxJe9uuWwA163HfZUCsfXXDA5IQeIFeSXvSu
d5/hq2mKYh0CkTqw27Dkt3yGY1sohoPI/mlKb3Ht1YktG3MTgN/GG8+HS2HB+danaemEM6uLM0fw
b7+9A6d0IG/mUCVehHMrG7t0Ohls+TF+uN0eSF4/YJp9xbDj0D8AUVddq7+cGLyPNmhHhwWdec+C
ThM9gjJmv36baRugTjpUJFY3FPm7zZUnM4/N2JX4yqBffiUM33U/QZzr7feIuOSMdEfd0/YYvBnJ
18NpRIrdSNC6ccqo1k+DE28hFQoHrC2E5MRSLaBOGrNMH2UCrEli5ME4irQ946rCaAXYvAZXJizF
+oBpn8qkUuHGzq7t3p9KBWoCpAeUBiaPfA/gps10IbMavMTvV9g9f06tk3e0Nqji44lAmRJIhe8U
76UPp2Px11gST40cBOJsJFTV5gTOx/MMHISaQtlBDRQeuXQySXQCqihm+QbrXwQ5KE4w888FnqjH
KlOGkozQr02tefMoYBzaAXa2gmx/kPCrffwaQ90TLiH8NLoYbaAoov8KcT+o6WtuaYcr1mFwIh6f
/KrJmiMXTkyTItAlR6KFoB4ORd87RMD3TWdj2eYsd5Ceyz+xQ6GbzpKtlQByfbzhtR/t7RrZ3rhd
mQ1pYEGUtEsMwlFNZAw4pLg6RO867dMc8Me/CEAA2d867RvRJcPIPBWLEmA+O/Axb7ojsaTmj6Ea
MALdJ04Gect6YpD/gE59QDKUrfrk3AJ1Jr2vFS04PIMFd09+YkiNAthSlW0m2Hw7Ar9S86D4Tmqd
NFSt1qd1Q4eKuQpaCdnCi4VTZa7y3iU0qImHBVyjpdH9LmkOFxSU3eeLnvC2smTCQ5ZSnJ0r06xB
4gdokT1Y13G1fMomZCRcF/wr7BC+VSib4bB91A2QkgeteJCA10OBpZNRY+ozOP8PaKUOmS+fcM4U
r4cqpwD4b7WmFXZec/FCNZ8xMFVgLihCNZEHGiQFjdaABRLue6eHZAoFSNEXf+okJ6CmUIn6MMa7
PxFcoTG4W97qI3Uy3S8WsRBDNwd6jndgVSt3c/TLYYWQCzENpIBnFD83dFob11UX2VOJrBCm78dr
vUGFgrf6+LqeV357b7qgqBDIUZdkJo7cbWWakD/DokMFb2YGgPnok9M5cH7WkNE/1gUgUTxcOA/O
p64+Vhy6ypZLecmzOMFgIEHUALvL3RowjtqrE7Oue8eT4rYpehMPmAxGlYIMPln5lO4IFfFt6ymP
C3x4ASoCXc2tRR4BOC92r+oPQu4NM52QXISk4BNqSdtoXSh54l4Vf/Zn1FiA95Y6pvg3Q63kLc4L
/jNyNFXwDimKw49oNay/4IrzFSZGTgmU9kdGB9Ov+7oloIg/E0sW4sgtjCxpzw75Bs3bRFJkAnLt
S29dO/mbyXFihzoU1XFzXbiNfj0bUGY73bZKercZ2+iNQBwphWjdOBDNMrSL4i+lg+F9TTzpAHmi
QndTFwLGclHmN2U20O33+b7UE/a06Aa7Q3OOyLKVTeez7IjiZNqIXtX+tryzsiWa4D9TLwIvr1mN
E2hoOSZk0RZxWVj7RQaFP56r5OUXMeEwtyqvmK6YDllb1IewDTSaqfeLw1+9b47bdujWb+rKwcUm
QzTIbHVgrXwgvoA21HYy87xl++t2wT1eDUGpWv67o4yff9FrSTs+D6uoGJqCemo2V2qqrdPMxZOv
r+PDDRkF6SVKMdz7F32TvAiRKmrZwMOKGYowTdonJ2ss2hrhc5z1Pj8vZ6xTVnQky8UfnSZteY5U
qYi/oWqb+TmbJIJcVL2Yjx4KXj7STQ3HZN3f9ke2sg81rzX5GnLmVTIWSGb0RPYCNS6zo5uAOvQe
mMXUsg77Qw5bnD93aZ7rApr7H90XS+8eVx4IN7PyPuZVgw1imxu2K+T1x3JMKQaTvjnrYA0vKVTI
HDT2Uh8PNzdO3oHVUFQCx+7qLewn9DOxz6PKTjKQQ029N5qnmmOH4rD13yJsgFY50woSiEzHVCov
tpBYUzpQGo/YZYdpI/adz6/MQbyvyoybaYUqpX/oNThBgVkrEN5Y5CKWfKjkJJSZhZZOEXH+beGJ
ZF2xCcam0Rbft7dSgo6NEE4RJLga353cBRY8DaN8bTuriMPPlk6/gIBuqTZ56x8eetzTx2v9fhZA
Sc1QUmNyQWbAAALI//CZNPwL8h9irIjwg9upIX4gxaZm8PhLPKB6Zr5YeWqZqGwqzwqMzPIlABQH
hnRBpXi1HOOjdjSgzhfW8VGcjdXMWQyCrK5dRbfGaOtXE3Ubm5h8LwIVYOTqU/YP61J4HzCw/2or
L/nRZmpaLUCQSi2D5BpbI3TXbP9mE8+Jj8UYuj18WvlWODs82phUvsn9t3vpf0aTlcCDSXgGndIx
S8rrq0ZBmRnHURRFBs0kghl8uFj/fUq+2RoWVhlhlF9ZbgyOlFOVEwtNpiWrgkRvVhmQPq6cfwcw
FgIFghhtRgNX90GEfE257EgNFyFE6kA6fDVTs5aq/AoExS9y7M3aeXRFSxwnMaa4fcodmfKM2QBy
Ui9CjYeJ+XDArKc/Sroa4MQ40E7rCHkvWUBgz8zYpeF05+uF2COT5YPZMITposcqyHWc7+etAt+Z
ZDN07t6kgxaiy3NgqIckBOIU7O2VwnQEqOALKtxR172CA2zk4+xkWHG5IQEc2TNavAinV/LaO7BP
ylYYDGb8M/aveqfHYgIMksnzSeRF2Q3AMnDt1BUD1LJZKJHdeuLWwetg9rCJARty2vjtgmL3Shap
kiVYOp/52sIe5ISgSuNoS6Qufiva3Acqimwfpeu5/qRs3QXp3mtr4SkpcHTPQfRmLKZW4EQGrhdv
z9xoP7aRDhcH2TvkOFyFnagfmVoaXZgihnGZzF8gg+5O+jtMgElRr8fLHOLuuF8zECZlslJXAlQK
2ujAvKunfvW0Iw0x9/zCeO1x4L0rT8LAk3IUn+tX3sct95hf7UAPt7X7gchwHuJzNtrB6/vGMVsY
swz7HzMwkG/kLgUc37B32BMKwgEYKMkTgPI2aLOgI3YiD+zLsFB7j3yyok6lFvNtpxUwi6IKgkuQ
YELAI9AEOIsjziadL6ntrdp0osb1wM+Yq0gSqlCocwkQ2ipOoC/79DpORJLIdvT9a3ELso1dFMi8
FlEsJCcgMlA/Nz20ZII7lfqj8GeVmwqZ7ZwbxwWSUodlfEMJWmeTEEAC//EzZFEE5zJ4Ec78r/GM
CBUxR4k2KM1ZpLKEHVrAWeRLRn+KFhzGzAAsLscCywrSnsPwv8wCZ78cODD4jZqB6UWrHAVxcUU9
ilu75GT1dbWU7wbguOum6xByaRgw1R0BGINJzzx55uwmdX5leVEhOZ1gF0fBjC1w3fqKoZfJi4ye
+/ix6ILXeSYPWTkuLGvz8SEYFbr7fKBv2OaIeX7qV+zZfzS0oHk1nBL2a47apR3u8ZdgDEi1F5Qy
O0b4ZNIkDcHp2V78Prfyfero+XI/jXcBu0EP9HQTpiLzdJYmnU6Wo/8ufwR16TfD8XnaySPx/cTC
3CqdGAdCWboZC/VJznMnAWv8DagdB7HDnA7P7TVTEeZyWY4xhycVVEB5W9CNdiSCBGt/U7s4eWs/
sOBi4R1q5zDRrcLp5bbPK39QC/v4v1hymQkuSK8YgDGeK/R/vdTpQmk78dmo/inWduggH3xGiHne
HdNaaQX5emctCxCEucr8ZZXwdTACTAIladvGn8wGN090z3i5ECEGYRNDLp+p4MsVpEqDWeXP72Ww
9sDDRzCQJM/lXOnMu91hW0aRMFcKhcCvRPbou9ZFyeXCAx9Srpd3Q9R+iVvfvLK45WheFLtVq5Yd
4l90NMJvlcFlhmjKpLANXl8kJ9LR0/NDfBU+rCnatzfHkhsDjMhD5agY0pslAVTtvAv+uJKXBI2G
2HWlnBJ3PP1dmLQ5beJ/tOoIUoeAc/nH2aU8TbL1wLvFTlBI1zmuOZxF0ERQCtQHxdzAUM/3fl4Q
/ukaHL+qQhn0r+Rn5CFNRcG4ah9jbSk/yR+uWym4f3mP9uS1+3e6EKgWsRCn1Tm+t83/xJWsgbY8
gc46j7XuUgC65GM1/euv/p4rP+BcTaVcEMT38Sw0/FDkgmmQii9eBLsx2lXhC3lhPgypc74v4bwE
3mkeQ/WODSBmHOkgLVvj0Y9TYqNKtJllsg8ejQekf/fIg3rHhCFkzBVfX9clNy4CAOEyCi6kFIvL
HRyiU+0JeAzgbShf82rOFiAPpEkOwOSDVk7K6BWRYuukfNuxibbg/KCrifE4oWZ+ipxDiyRCnyKI
uRGOKxKiK8uk4Dmf2YNGA+bUDXqLkwHCe6o4OSGYf6BdtdTrsEbPqudANAzFt+sQOZB65aD2cQZN
n83Vgn/lbJ95EeMSHyhoiJLCr3csXMCwT6ivUiUQ8e/kzawIkZk2dr0ZDOerusaSXuh6XoRmuN5x
RyPVoWAHkGkXWt70iVLPXfBwd8UJ7R2g2EfdDBUivSK0+ly/+SlkZ9scrhDBqq9LwjD0PhlYYYpu
a5L5tkxqxz0tX3HQ4GzhNifBf2T3lD4wGrD9jPNrJ41o8E8BWQ9lCXQqg2OM3cLJe+Vdkq2rAuMq
zwAcEOMvgnpuTid5venvWbCk0FZoQr9VA4RoxiLY6ABKjI7u4S80r7XtNrjNBLYzOb5/Vk6ODxdO
jCDheXSckNVSA5R5AwTpxl4mtN8stL4MzsyQafZcrimbTnwxbBZS5B652NsneG92JBHJLFCGv95t
SWHRbIIVQTB+xAXihnUXga7lYMy1t+Gbc/d6Vg5L1iLhIXX2vVhvyvXA56axaTWPAuu1LbzzlHkD
WhNv+ucWfIrk9SqBshQWmMkzBK0o5N+4Goyo+/OIyUgETDfCUmIaXLUQ8rU8F4cvPRLnl/s8hL3B
fxheAkOy8piW0mU4wR93PG7qU/qwesInnF/7ozTKzYvKptinup1rQfMevm8f+HXlov2J0rx/HmQr
t5LK/Yd/t5sm+ryTubHxfmh79OULAqTJl2IaN/8lrFm/4b7prFwwptU8z95E94ML/6LC2Pe8X8Q2
pWZEEHkg0g9xYlB3DFx7q4BcIvuQKOHf52jeYRi2lYuebcEaFBiOaPfR+hcao9+81u049j2A8TMo
4BV7xc/OH5/AiUoMM80S6wwmfKMEOCjb6AI810+CzKoEk1OCSL5G1DIc+uKfWLAzuE0yQJOoe4Tl
mx4b8DAvZuTeand/JT+4gLK/wzcP18Mv/O+HMSDFFjWG7QbxTa2Wf+umSmfi5UAzMiCP1g81te+S
o/ritKMzCPDQ71MgHdBmzbPNb+rW+rZzNe66eHyAypcTRy0sRx10YNkaL0TklY8DAqC9+DxgI2dG
Pt1vuX/brXTHtzZoniu9EnRMxS93gjfFwE+2tjSny1wgNfNWJ19C6stY+xPJsXHq+Xkx11XBXjkM
kRlvRHrmyIBW49YySlOpXu1BRAFmHpLbxauEUVk0HoLDMQjiDUiUneQVVTFpkC37CqpDJYxdqd0f
TB6tz9/GyTzkvKBjcQf5CUF58MJDn8RXiZrsHHy2JsC9gCtpeKTcl6WIHJnG9oUrcK13zka1aC7r
2TwS2AN6Iv6etbJRVJy6EufTAAlICXFNTdbVphoYoOpPmWNuG0YvccYSHbnVecrlXzzQIIMkP+ea
YgsT4SOeLG1WUBEw1PmEU9XOK1HcF734hxdZ0QPFM7CDSE6AzKerTs/kcUvKyYsjWG281HkU4cRp
DigLbRXjgM2LIZPTBH2v7ihrLEDyLTkUNYBzgsnI6omh1cBgVptoCWAS39cVE5cruceh5NRL3M+E
aRovSbi2W9//iKScolIC7GjmyA4WF52POf2h0yan471rMCHiWsrEzqbMJoQwu9Clac7u5+3vOmiu
kjO+La1sY28h2VbKDTUFfBBxSI8bxw/pjpeFY9zWVkIphT5FYvAkx2YFiSxPQ/A7/hu2/kSRBGBV
xUoCm2tW9hZ5xZakVn2DEYF1ikjmx5MauiUmGCQoeJPxSkAxpt4k+7u/JZeejP09/m+m76G8uJ0c
4gXBCjGnhQWizJSsBAkjKAQxPCEKl/A7wPVZ5Nh/LMKciYqetFPPv1nJNjEODfVGn06t5HhVpuAE
O1Pxb1apv7DBHTNcGjzQlCLIBgPSVD/gxhFFoc+rfcG6yPG94z0G6B0ldIr4583bVce6b7b7uHMe
AxMoVkecBICKuI//mbaAOKRhUSx3NBxWDiS1zSW6DEHYN77hFn8l3XBEPVPhzi20zdnM8xfTTjpB
PrCTYscsgE92O2/XM3XlDeisvYIvcirRjghO92tdGlo0DA3O+F+RcUHJTkUn4y0IG4e4FDycCCdr
Qzfwpt//3f57irT79JqYNUEmDbDx/pkVYZCSHsUaXBeWWEOfj0wOouVBkCH+qfVAqtFbxslouIA9
P8QGgu639ol0oG0kLzn4scTut11jm55BFvS5b/cMpR480stzoj0smyDrwKs2OGcjohIUMsP8RlPq
Un1NZGfcEmx/EdLXM9gToSIQJcWlfxLN1K1rK/VJ3+pQt1QqFdyGL3G8vUFuvPAtoh2gdu9uaVDx
YvRoV4AsXbO54hClmjVLyUtufeiMjoL14ankkI/I9MSPGmMfBSreBkIJDt2tMbniYYcQ6HEsXGU+
ha7KJj6TETqx2RSvxOFHcVJPOlLPZkWP+xG6MnBs7qsCd0ZB1bVkzrB31z0KJ7QpYfeZfEodUkbC
zWj+01djyE5pE+hqrr2JhisOe5BVwtRDuTejtrQJPmIqM9decsgWPVMHUVRWuQ+hb76XOuTsfrie
EZGzPw1VoB6mvAH39nXHLUM3BbUR0u+M47fvtWTN1oTC6ZKEwt/zo9ln79XZeMdchtdavxzGgyD7
OxUBBEGMtthZgQ2dQorJSx4DLQ8atnrqXUihsIIv67Csi2WQrOKRekLOncYrHhOaj7+3BpwYu7en
+Qc0aQYTIaWM6G8C3K8AyFd21s8TRcU271OG6Tb/Xr6UoW+a5jp5kMKnIvM8LjGNpoGoZwGdFhwU
ZgAuqcD3wcwZCG2czfETcgm1sX+jVbJSb+e+xJe+HUNtwJ6AIahtNrvp4Wr+7KQQ84wH3LBv7/0S
LbMq+LqNt4KnaD6nG6xvyyhUpN5SshmYNM6URlqQ25clNHkitokneHtiVriu+mFP6VAEEj3vPGTg
+9oT0XuIedq6sxN360Etjp/yAiGuDAYwL6yqqEv2vuZcevwTBrkA2fAbR3/ax7iASMc84r31pLd2
f4ykeBuYiraO4fBebyRDp/i7z3JPCXj934pQuV1WVjK5O4dhF4F5oU5qEbbzc3v5rrAbH7Wsqezt
KQhUsPAWkDV2cuwKjWTHq9lEARAdpr2ih5BpYyCwWvYCWpOXEi6NCqy++N+uoEHKo7pHhSKDqicX
057UynR02lAXX0CAN9lGZfkyW8WO6wSPcnJFrVZqBR3jpe2oyxcbV8nYrpA5sX14/WvaxmhR3RBi
+StC0d++7mqVa4ldJpJ6RY8wuWT5Ah4Is3NntvJTBu3dx0yarv6lLfGApiUNAobxmIFa9XTh4si/
kpZkkclhzMyGzSYrTIxbi6+sZDclTseOdve1lWik/pJnL5wIYjuRiPdt1+1WsIblT9C2TM1OUDi2
dINpbDqhmzxtobtBQVfYUjDTPDAO39IBYGFhXDN5DesgESfFkfoW5xGaNjFPfncl8PF7+rBap82n
KsJPtA938cvOudHwwUzafaPo3vqOCu/yrvZtc3SKklFCzPz1Ai/5RgdkQJMRk3v/Va4M4yBAF9Vj
7//sUYfs0Zgoe//Qri4VoTx+OLkZZBQE8JJcF4zsbvp6uGv9GZYrX+GmjbN7dCzLTY29a7tKam9o
3NfizkGagZQtZUveyt4E/NaClSvOKFHNO2jGPrHv00jdStbEgyGZa23KRn1lqUCxnTE9IdvGf6cT
LFcsZwozYTjxVleAOTMeX56wIkqsIjy8Hyl1ukmxoSDsyi8/l2iDhmPPiXfPGMSu/92etNXWlnph
fs7wLv0fwlhgvGfM6lMaZQ/zqI3iwBbh/55XhDYgsTe/vPCh2j3dh4DhSajPIwmn0qw8xxWB8IHD
HLxZPq7lIKVsEq0kau3/p76ZlZm/+2lPVo2P1xENVw93S1BAXFyVCBpsi+AAIgCH5Cby8YSKvqUo
dT2W/cK7TENfTmHiPcX/1Wx+nTs65l/FN3TWJNO0Pz0uk+IMoYr3BU859+9Ht2Wf6ciVJBySmahT
sNHo2nT9e0v5YB8f3zLi7pX6aZgMBA/YjkIhk1zI6aqwgvT2zBMeEVmEiWXkEn9Hc/mEj0mB73v8
9d7ptnqg2N2Ozl2c9muG+zaG/cZoiP1JyB1Qol+/d2FH+m80XrCbm/vpMszz/dsnlnmu2G7FUHQ+
mJd+59ecM2ny5rtbQISygQAeDWTtnkaZnoGuZ18cqCfxf2U5XGHkoN/ssRSKZW1+qrIGDF82CCgu
a9mDf9e6o3Z7TPCs6x+YAr+eoGplrCE9umGdnuYft6ZhYFsJs7ZH60UOXS4xNCzIXajxs44oj5+h
wiaT8w/9etcLUgwmf5LBQEkKQmEBw8Rcle8U8W9QNtZN4xN9VKJPzomje0L447pK4efTRt+sbjcp
N/x+Z+GB6O8XmBlr9HSgkoA77IxTsowDI/54vjmVxF3t1sb4tD6u1ksayIObXRFEwfOVWalPh8D8
68lt228cZZirebomX9RK0Ds52f6yDaWxs7mDzm1craMNs1S0J7UIQ6CP0qvVXd/vstNUy3C/K2Zp
fwjujOGkKbB5Y7UeXTEK+0pyDjxNVyfhIQrUUkcFch1r5T4kxrhfEAGQOJK60//9XN1HBvMxthLW
yNe/XvasK2Zq6mrmyirzAtjYP7wb+u8daWHzs1Ab1kQuxcgMwxjx+PRGF8Ndmf4JNj3sxQt/kunx
OeOg5RCp/TzV73Li4+e4qanDPrObHCq4Sbh1rwvUr+Xh6P7YzbbsT27spKCwA4mjC63y29fo32+Z
cUHYhD+29VFTlcFMZRpdXCOeepfdNZZOrW5xfITaN4xcug+bHgSTZvBu6x5+pHVadVTYRPl5rymC
ihKdEjTzza8dTNak0VU/PgnaEm68QtsxiZljj1ZLv601y68Q8/35n7ksDOU8eRPVZ8vue5Yqsyyd
CruJ4jN/BcubNax5XNmm4okUWyAoR47gLwmzPfC3IZNJ7tPNvI5cGkBYHLeP+h0hguIAgfNQYzqF
6DrmFAuVMZFLRmz2nDcpIZ6jr9JvIMf+yij/JCK0VF8VTUIT0gEbzJHAFFH7wCvFpWl31fZ+yl5K
F4DJGBusqEEQjjfpf0HG75xFVVfJLoy34AFG73muZcjac425BWUdWu+Kfw1D9bZdsyujI7sqGJ8z
epBZ7uX78SFRRYGLVCmqNNO7GFnf8E9PeSNvSlUKmab0VaEsiGpPVtmewNDM5fRKog3WrP/VwJa8
LzyHy/JnvPSVLOM2eFe8Z5pafR7L0uwIYUEnLuUe/YU4pwao8vbdOjGmF8pWYPH4wlqRq+xzzMOq
tKdHN+VX2vMXnHF66jxeGbkaCL+SgcDevKYGSmrHi7KVN6v3xPTV3f0GUq9F1fkheN5M9ProVKtu
rhovj6rDEVenwVLiLISt/1zwCsZSK7qal4ygbmpOKBr6VMykJy2YNA9XKLQUtHYwj4FAVQHLv3s5
Qy+P2Dd7c5EpXaQYIW89YJMPB8kT9e84D1Tv/LK05dcZ6u4kzFhZH8w55fqrjnRrEH1EQIigDxxc
4cAOGr6vW0g0GISUxxN8JzI9KvXsLRpLRqHIichzxBdz+UTUR+A+KG2+n5Y1yb+CUr9EgdbqDXa7
xeIJtRMO1T7j1ouV7vUHfW70M+OpiJ35JFTNEB+AKVBJGGAoGjA59m1EEiXSVwEY/owIgfK2vwwf
QisLbdg9Qu0PQI4lU2g+DSvxr4ylyF8IcOsvVA3iWtNTLJrnRPT/6PKxBCpgamxaGSwmsfE7tcwO
7Yw6thEZMs2gYzak8BodwJVvanuNFm2MTb7UDdbvRyquwoZob+hhPnCnsofAvVfl7xMqzWUwREm+
Y8/6Tvoww9OD38UzNAtknliSjY6e++3f1jHAKRE8zFLSlaJujc71qrVEOzRDRfosA3BEhYSy3Mbm
9qR/imTJRA3V7lwtUxqOqaRWuBuadOvhrjDGOLxvultcgBGqAmkwC35IbKsiaB6bqQZxweAyE/1Y
dBs7Z6rkk+MOU2kIHIEsQCGiivUd9ltfPsLykv02Lu4VFtYd9P3TI8Ct3V0d5qhXSQUPAb3dhuOP
Gt08BSK/bS6hoEyUqylUBYqBlrqYC359pE2TSeMhfRCG/YYulPCS2xGdCs3C4xHQjtduhGRX5XHG
FrPIiaf5OnUcBhcdvO2fJuCtvJDYlqBjmznGzk8KzGp3nGFzMtbCmEm2P1r5twHJvwaf2QN2NR+4
361MEFlelsrwyBgY7FVxB1iks0cNZCUUbPkrsDX/2v9ZyNtuKX2PfJFjHCBbcikpGNIWae7pPvvV
yPdW1Ei1/eDBifiBdfQDqJS1wo4s7sufTIsl2lAuLso4F4mTOwSSyfhvpGacdV53EKr3MP1DxAeI
mfvWEZ4i0dm4Au52Gai4apWZ00DXe0XYAFK51ottkpoKN6Ew+fT2Uxyn6uKCqVgOlSwU7oKPnqYS
2E7KmmkEtc269zXKYtW7iYf3ePiSo1s1nXSPf49Roo8rvouyGblI9rwH+4WmJEIknKgqW4l/sa3y
Tgv0AuTvCBfcTm4hQ9+0uxcj/Zd0p5QMesSueB3sHiXZdjGUO9lSVFUbq/VS+t7ABLVVvYzHJMyQ
T9utg1SSAGCkPogZXv9atQrwQnuvak13KVFYHGDLu0zk5Xlhd8hnBTxXZVyh8vf/w1h6ZooEzGg3
9KSS0v/e6eLIlcxZJveqEW2X/7AdD04699WuMAkxqFNDDlp0Ivrwz6kxFFtKBmIdAkIWXciBzu1h
uEeMi/jvDnHnYUZZHumEetQBadt3whe6zT58c2ufMyxO41UsRgCBFtC/ZzLNCIambwdq0ZoAr75H
YXcNX3Ws681rxnhS3GkAhQUhMSNj90Cx6UJ8AXMS/QmPptK2osnIEH2dcwC1pDBZ+Ovi5nlDSTnF
7xLqP4N36k5x6VMW59AS7QKZTzQAkkhujZhvbLLHTQyxrNCrIhT2rc+F+x5IvjGxpu7LB2XSsGVS
GHVj3GUKwpRQWDdTWCOpE4Ob/Rd83Emh5+nmDWaz7SOf00+jzf6TCnQDiG3TOwr5wifhRo+zNa7w
834cegRdOv0q46YQGAEMC/C3TNmrhuuiVE3KOqDhMsXVg8bVKK1K9MOYl0xSDc+8sa3CmWGJvDp/
ZywgtuwaZUEuN7C1ZFj0mIL//UCuHGicY0gjL1mRqMqGwsgQ/fwk5F3eMBwa/XGD6mEbEfjetH3S
BRiB8GcHF/oy5NoakMPFdtTgKWCxxk7h1KQdZ/q6A3u+EhWd5Lm6moGiarzIPKlCibTAsfe7i7B/
4SerCEMXzwlpi9sb09iNsRcoavQaNeX1o4dN4/8UqRxrAXgTL23tIE6FyeT8dKT4RmLjr+kX+jmh
A0u9a1nBp6AJU4EeRkRnV7MRj3c678pJicMVLZVGISMSwuoW/4FikviGnwQTQXkgD6n0VLjqIN5l
ta2e7vtl/vuwhYYvUbXQW0EGPorHrhod/dljl1uWijDFFloMCZZY+zxKtWtd4grWwUpIuPUBeOkK
yZfieYaJv43/l8/zMVnDRDNw7qTVp3+A36fJBZJaepBCMkeCUMe2WXIc2rzfvAYBshRVlOUR3kPL
AI3GKxVQXjIjZbhb7eFH5rpojImx7BFHfl+9MDBbP8KRqSJLDinr8QvZJOX3E/anxvTsqb41Gtgd
Ru9TKHq+96HKw+kL7A7OH+/Cj4eRCy3+YOWeUASlXffp6FqClLq3HwTQ3Be39bq1ffLKVLXqbuhi
ffV62rbWSd6bqRnzYsrw/WqQybPJP6akA8kGKOvwj9oJNb0PAIKZfeWZSZ+Eq6W6cqP4llub6/H9
KsKKY9Op/J+ML+NMC+oshCka/q8MI6JStSljMW5Jlz55b66TtPUiE2SzsPTEvsSuYvMdr44eJsDo
g0eLNDU6IF359xx/C39JUKUXZ9IFSjk1dd7isXNijfOsectk8jkXfTPH7/EV7/r7LJrRjRgJq0+/
qolRbqjSAFxXEWk2qPhfhO4wAF4ebgqy8yeP7JEb9NA1Cwua0Z0uewta4UBnZb5CYuc39qjq35/r
nFK4zlRR3WuPuwThpRwWC9a2M4qcYniNEIFhM1LvjjbViRHmReuCbB1YjAaCvOfT/cHEYwlq6dIr
J0OF0/oNKJ0Loil/pz2ZxgMBvxSHwtXMfkdO7dImeSZMlO30inTJXNZcS5wZBVFErQNl41v6rV22
VG49GZmw9qt90MoLozE+4x9Uezpl5ISCgSGGAq3yNcRxywPJdf7KmLIKqki8AhrOX70K/LGS2o5A
/iZvAUowIUea/nNkFf/WJwl+JY52LXo8f6T2DzAzAkLjuLHdHrlfbfaUwSpkwehmkGPZbb4nFoVV
tZKbDWRWxHuHKORvR1YXLt9iG1jGd3ai/lkJzoca3mAmmklzFaN4kxR9K9LpJZSjtwM680g4LsVS
HDDFnTJV1iqBrnn9z888siy89z3xqmU2Vtbf9lBM5ZAFKybTNKSGhXFy8oEfSpxDiQBwbT4X82/g
4CkqN0QIeMx3t3j+AgFAwGa2AYStMCuEhrz4LDtnfyt0uSI+6E/hrZ0Mw8PCc/lU1aa8dCT0d7YW
bn5QQvIrVomOCGNIXNsEeIJmBvdBUDj5McvCevO1vXzyPSBRermSxI5Od46EehyDXRU4bwfeY0Si
HjOYWb/2N6e23tQGHL0A03zfgA7E7p2xydI1zKRYmBzMwRcI5f7vATSgAtCi58c6ZO+SvT1LUhmK
IcQKBW059XtRXVCV654sSCjB/TlPw+ylZ35u1Wffb+B0a35BZgFqQ/9IHhtfSYV35pOSOyUI0yz5
jd2Q596O8vRDSZhlKecgUbUPdPMvcqdihl3RudtlWk3YDF+W7BZWKY8uk+nOp9EnSkQidf1Sr8BC
FT9yoEuj8tW3sfD3y6peoDxjLODeDmZKDaJQmvbr09vnHlvleYX9Ia2HST32AN7lTq+ZHBcJGa/O
+ww46kb2KafQIRPd7ZvN/jOG2Ozc2r+6ruEctLM7jocp1AtQwnWdgW8T1P387oM3/whMRO8ieq8p
Muzt3ufkem9kCCxQdrhdTlcj3CkkTZmIdnoPAOja/UOZGzAMqdZV85dRK8Q5Z98j20ULAb6pmK2T
u3pRWErv5jlKbqvswjj1egO2lBSb8tfRlGNUrSvgeUkvwL1to3P1Er0WF2vXvELx9sqeF3V3oYal
dG3ec5Wu2SZ33//kfCfTp8hDyEyHDkQicSDnd3/XwohBHpyZRiuwCbuNpeUzBGDuPMDNtgRFL0qp
qU9fwRvFaNqgSlBwIaAs4smDzHqXg0h4SkyPLOC7iglcxdjUzXfFQ2J237YStDEi2F5cghAhxxFE
arxzAkOkdj0ScZbmiKY6sykQ2VfL++ekm0KYtv8341XmVvN1o8UnoTYjZOYMOPj3BgX/XE9oag5S
ul4z1Sy7yQL4HUbzNkTmBS81hFOroVyNbliZ+wsW2fjZpHKvABZ/bwOATer/lb+TaCSRLRERnLmT
4yOynqFKK9FIPVCmaOik93FOg52ZiK6yHGkJm5dC1SrC3cf9pk8/PUL8bi+EbsVinWl9RHfy1LXH
64fz3PIQXnfAUxpankvYhBJ60E59JzMFiIOJwsYkFuWcDoNwUkw0qEN1SRag3ibbZcbdeq6mYV+U
OXzPTlHyTpKZpn+rVxN96PrOmEMN/4GvQUrkGwkL6PlOCvLHjrcQrn9P6PrvfxqFjVfm4tz0HQtJ
WIF/ui0MhsSMLPd70pVZS34hIKMemfPdhs/EbZxigu1dIzNcen91hx+b9aPpRzmW3j8cUlgXKDrq
2Skt8kTXvkEXhwIJHlNi04y8SqYJY6ccXb8EMK/Kau/CfQa4AeMzfvx6cNKTDlAN5eZCZKGS5Loh
oA3+mxJLXDcrpwpDKNrur3R1iMqngWwEoBFqtXlfaMEN1RtCOEoUCuTLxk6LA0SO54ssd8B31XVF
83fQpd/YW26MyW7tjbfi8WID6ERFVGVGEmQMxAvxKfz2Ulc33lyZB2A3o4nvZN+cHVAOY2ScGokQ
CtrDwhXljRZ3/xdSRogQJFZ5o84LZbgx9e5WVgnPvLj9ammF4H+RRt6EL/Rb0uSFESao9rxRseBU
Qjy4M2so++EAHXCTUQqombeCZRjH4chb9tbu31EU7BWwwqLTxiR44vwaH/w3+2wlfKwaYHKb2/Y3
gXeMB3ksrfSHVjn21TkYfj1CJRmDBMMlcmCCM0URJNbTaikpesYX5ZlaCNgSZhfecp32Fublu8bl
h24gPAdfgM523WbPoyzwlUHi5haFlmuKpJyYqbJtMSrvvI5p0OOBBuWV1H0+UrJ2PO1pTpRv4K4Q
TO9CePoN5eMs9n6aF4cYwrR7Q+hsnaawo2AAyvPsCcTuO4npnadvps/YM+9ihpGeGeQnhlhnvzew
OofkV/Eqqcdo6bs5akhunAOLnUo1oaY6y2s3U3HQsYhA5T49ALXyvzeVso9CcrMpmIhc2aqkxYR6
3t/4NrzC47KvE9j9Jew0I00TxKOUYiU51LwVLrqPVi19rRuL5B74CozEULmG+i2DCbbnlzNBu8oR
xfRTGO3nKAfIajQX92hEvFzmiN4UFTe/DBbwOAsmHsvfrFIITGza+CQbo536KhGmacV7tfHWjKji
hfarRKs1ZI8Ygz6xYQm8QIXYuh8D0CQEhw1TvkvZOANP4AfVihmM4kAp3jY/yJI03Zg770e/qm1i
CxIR99DU6C2YV4F8otMu5lqIRn5xB9g4PMxjb5BP7XSCnEWbqrf/i/6CcjBLYmLsNk5Ncbc05B7S
KnHM1L/UEbZLmK0ht0/vl+8wL8dGowz2LzlFIPAB5OuUjKJzYxb+3s9T0w+2fQ9IWt3+KWiXdbmK
/MUR9LKdCxFR6t780hBKJQpGzYXNSSiKg8BTS2BzwDC4KIb0+l+Owe4YEJACRE1GWFAs4N4YNKD/
UFPSnm3Tjfze18Vrx4ZSCxHzXwSP11MlOg9bybSGOZBTKPh0j31PNjlQyd7GJK2oKrD5JuaAxLRU
uHahH+NaikNnkwAyZGquDSGIPwBlCrdm5gih2kunVoLgCxkGuX2H1ylrxJmKrW08tMcC0nRvjFUH
tDTm5NhE0QVhXdEKOq9GIi9iZD/tIsGOWf43/lo3nMR9sccPHs74esgoDEXCtA4YouNFslPnhUEc
zYhDbGmqCIE4rMreHpuZnfSSHmFnp9wMBncQWALtJJ1hTQUiVJ7gRXibLMSJEMxXbyyn2EJTczE3
NDD3GfHsuxvQMB2YOUneBdlna1PMROYCN8RfsDNmibDqftECgCsrt84boYG05Srv0CdlNWayxJs2
k3G9LNlwG2Equ6a9nfeddfUrFcZPiFGFjDd9DK7RU3R0RQA9Y1xlAYSfxqi9DsReMeAgedOQ773+
ywKhp+oS2pAACzJqIwAp5hWAPy951UVL6IwZo2Wjj6EdJ+ZEe4RFidFcfDyVNFgbTiCNOncrFmcd
dARgVxsQDI7eRxMCWEmHwKjeI4j2N/Xp56pmiPyjtnevP7ndbN7WTEW9kuTqy+rsie/qgyH8fYDI
fRzvo3SNghtF3y57OB9CCfIQPSLvvMaYGUCDKwzD4s8JMprhf6bMSgIf5FIa9b4NcZDQv8E1ln50
yzgvvNSV9yxmQjUacvyaQgx8KHQ+wcGmd+QvHRokkgy+qGleE6mIppJdxNc8O2hPofWjy7AVdKZu
usr/atVl7WwJ2UTEN4vosA439nyw7bxJn6NaaociKpHqTs7RDFU87VIHIzDUPBAWpBtx0r0iCzgP
MCelcp5WFk9GgN3nNC0sycP8DqUdddra6cYlR1PGhLI6WKA6Zg4IQTv8K7gff/yNjF/m97Bgwqcw
y8T4Fit6DqDZeQD/snoQuMWXVTUVFehjoHGE8do2ajfoCwHn12L4OY2ugr9++8poGSvsnNd7BW/T
IHs4jvHWJD/vILRY0h5yPOT2gwDy1cHO/vniReo4Cb6uwFYyJoupwj/ASW1AaNyvesws1lkvH00d
Rn6tF5NTRnwJrSaiWs5t4WI6icyltjkGKgXgMJPZsp5CQloYSPJfOAIiNud4iJEOygC06K6xv9w8
kYvDnQwDW2moGloS37PLo6qI916l/yxFBYeHSoHXqWErtGGRrjo/ntwxGV86C/9oPEYnXZzqGmF1
OHRiE1qC3guX/odN0C25m54zKnFtj3u/dsfrA9jsKotQxd+RX5xZr4fy0JGmorQm5gmO4bd8Wda+
cbIBUwKhPQy9HMMAXoWuaDQdXcug2ko6lFaExUySaf1HKH0NVhNExjV4sWzhw1YRZ4q0BSbgB//m
U/rsvGmUJSSLsBZtg6VSICMsoa+e8pnLKVT0Mfrhv8HQ8YVlF5U+AFd2BBM/p1UopxqEg5+jUrd5
/rdEFv4dwiA5osHjRXImA0vHP0N6H+pLIfB1EzZRaNad16OCi62q0ljNZVXy0WRgofsY6gyaudQD
iP2Uw02cEsQYIZFoWCF6JHrkgEzag8l2b+C5b5q1nn4ko4btv7cpvs89Ke/3mvJoKZ2zpmVoHJfu
NPKiJ3Qt1OZNgvW17dyJQtoeTSWkfJ1GbItt7j5wUHXYcUk3QVLq6b6AeVKizm4ivKOZ9X7ZSnBS
VVB40utWReq7/8NgD1Q8dkQZf1H32L2U/wtbTK3eGEsao5AZ1+Dlf82Ra9aAlMghQx3za/jT4j6z
zL3xELH4rNl4AZ7EKMJnyWgweubvfFOa/Wh1Y8erLFjufg8K6W79E0uA1A4QxxgVNcR5lqS1obj1
E4jv8gFVx0AfrkonIJh/44D/rskS8IUxFN+xLihhdjmpK2zLntaWD4Q40VST5CFlHcQFEm144kxZ
4ztmU9QLTL01kxpUQsKgTy3HolhxNW1lLLwAlLdNcFDrm5FEZKu/wv7pd25iFJFJ/7AwoCIMzZc0
mLpi5rFYdL0nyPJWcogWNWGLMmuCpa3DlODX7/LlQnEUeJEvY4+TnbryuGbjF4mwToRRYl2X/sT0
iTsCxKkECN8Eep766EXvy+oImXQ+PxzGukRNojGT+mMAOpWQvIJ6Gzd8lCHeLrorJK3UavPYq3pd
icKrS8PV/VGb9O42Bf4BxiEvm9MRMgXlPInVdIGSKYwAt+Y96tGncE4PjaIBynVL43pz+B2rHmZa
uXbkt44IxXpkzxD5JAf6BTj8M87v3JnHupubcNVLfyRbs4FdMqPDcjwzEaFyVUbwjqx9rxSE6Ogg
rM//gCJjxGTzdWgD9tsLe7U3eSOIdbvh1HRwMXJjRFmo2GU6Y4k+93eXV+MBYdwnMnd9Oey1G2dz
be0do+XCg1JSNZ0RzIG2FsLfSV0/T2FLaOYrikSh+77g+4VgoZnWv/c2hD1V0SGGvzUf2sWBO8GN
3UQB/xONlJ2O6UYiOkjUKLoTqsKAruDWBO5IPdg4BB2mqIJn5h26q6XACyK2y3IdPM+U4Lxt9d5K
5MoAtXfMG+g2ljxf6xSULR7m7ObIqUPOcJcwtmIst85ntkXb7Uc1EezJFJ5rVrwEz6Nq4CnXGxIX
t2SJBeHnq0qqnOiEJE1vJ60nRN0xLYtRitm+Rk3By1fkTlF74DP1MmHUCR4owRDAHa/jBzz4oK20
CVzNrH6oA10HpHtNNnY8zLwXqeCfnG0cv1bVCoFM4qIKB+1p5J25CSjjsh2iI9G6t2Jgvh+ZBUdf
WbSVyfozooVeaty8A5ZmoTEf2WaNvnCyOT4M5A/EvLwJ+akCG2Rx/xtB6wj7BJam97GaTwWmekh6
7nzep8Ocv5QC4NKYKQTlyrpEXIy6zTmem+sgBqMYMUqg9LIRp8c8lHt6uOseRXe9sp3wyXpAav7K
cjRyjBN8x1f56DbR1xXYQIFYYQO2Fwmjhtko/r4babeXwqln+yRg2A439pH8xKeNdYxWtOscyEfJ
g10Qh22eSUK+W4VmCMzm9maGzzYxTO2eGvBLuZxfWM5JijIDdiGXx5W6FM62cvXRKAQGiK62pYyq
Rgg7oNUb85L/PzZgVbFsb1ZzjxlLjRf+XbcGyWiuGTP+Q1fvpJn43/2FSx+WHOmcCQyX9cLLsmd5
bcg3qN9y2IA23Zyu+CnCBxvfkicC3LciGEydGtlJuDJJCfXfNOVcQI9cq/BWDZs7cdjeCsePClk1
VDyVZ4QXybpkr1Kjt3zo4o9ssNBhce+bWt/r7Mn1Dm2NAvMfa72aQ5+d0xFr2OHPi0t9WsHNooGS
p4XbDcL1Hl96tAz+K9IJR/dUcjTA28+YR/hUIDfM/ycr1hkPO0+hPrdCm6uIb6YiAZCRW6+4Ughh
Q78gKlxLXp1isYDoOnX8qRAkgSLYX1GDmDom/0JSvaejANMaY/h6+ArvFKpzT4Lfignztv6xCiCu
IAgA8M7bwk3NcLGo95dWOFiIYe9sgSRI9gk5AhrnZPx+cqFlOfLkDiqTORll4pA7oKxq6xfuqJv4
QGTQPCfLnxsOWz+HH/S0e60gvDvWIsJ7GATEoD+s3bswynrMwiBXc3OlOj75mEqm+xF75gkMwcUB
DYDZBeSUg6ffFd8joWiVkGlwEyNkkrMQ+qVFPM+LAoOA8DL+Txj+njzrj4V+j2YBdTsIxkxYE64y
WW8hpEVoxpn8ve8kKlSFC+fiP0tHcwceascnk/6a9oBIkoVeo70xfOJT1ajo4iTmPF91M+7doUnM
TyxPsC6ckIHlts0PdQ3YB3x4Ga9UvIOT4gJ82YqryjAOtEn1VetB7yiHdzLl/5D4oSER7WNHNOFp
slnPLXO7Ks/ioNpiLefLFGV8g9Dv+c3JpMjZsfH53p+yTdDWp/S0cUfoiuwqBFjJLM08ZfLFf1u8
MnsuIcClkZzsG51FROLmzQXjn7xQCZjJmtOkR99sbQBEhT6tzL2GwO8MyeljEvGAfnYB7XsDTmIU
h8brn4YSCga8cyF5XYLp+S54nhfn79dYLF/CvlR31Z/xCWJsiSEt6kFktUyBs35Gy+QRBYxwknOV
QtJIyoKRp1S9184aM4p1aXOok36Jv4iOiJIE7sxKOWKgNcJq6GCy+zhrh99szeKAtifOiZTmtNGM
aq3USoQ+O5I/XxqxgBakmJb6Cze4vZM9mTBqJo8SvSTfBzo2LyXxrytpppdFI+yb4IHiZR+LMvvr
3F333zw69HW6jIKhaYdmzmT45uH3zcdFBoY5mB0kWEld0b3XgSfBGfZ6GVSa3W92pLEs5rj4lTtb
T64lli4nqcO9nouvTngeaXeO05nmMK6eW7RV+mhPuCzhtW81jQKr+DUrmTJJg+rsM3wWDNEGereK
WuIFr44ClYYicgyoZk5lDHyGJueMm+kmVSGsN2pwE8MNq/8Vo8CzGmNQfRKT3dOfyecfTVnQQd6P
qMjS3Jaa01UiwGtW9oV8WPZBNU8gIplJ6QhCcvxgS2zpRGGsd2oSM2bNOW0iZ6dOr8d5bi7kkspi
OIm8rhUM0u/Xg62BwPGqIT9o7shuK3r9KzvjCDqML+2hU9SZPvOcsA9/25fyv2F+ertTDcoVVm+0
/ULi3hY5TEjKaD0QQ7fvPX7NjR2O7uOetdIZYFZNjhlFUEL/ukiVjAtZDVwBuKBUKiLMizxiS1zx
3lD1VsQY29iGzgDQ3kYrXa9rLnFo5C21cughtbeTLC76epwfCEXBaKepxQ9vS313NDsY55ddQpZn
nRA/cX2L5PD0bsiGv9xWm54fFBo7V6F5zNrcf80bChCaviDYr2UC4DQQg+VrnP59tEsH+rdmDYWy
/9/7aMzMwn4+jGtcNH3XoPAlgasyLwoZSqXQ58aQPkiFDejEWNT4PqB+FEHTSUtP1bIniTpttQuD
jzzZX5h7pcOBcR6JPftXmvNYzWBZWTRb5Uvtq/LDu6CX1gpKAcXe876Ll9B1ntTbetH+8qm+1gHx
ueHtVt6pzoy6CfUMXHvV7akA8dPndknuvJqwW+tYMmK6tkVA84ElztFn0fQepVNApTFATc6AHBev
dx93Vb6A0z3+CmYFH55tmeqemevuhJ+/UEyn/QzGWeAuM3wkkr8pcxmx6S3wa37DoXzCvjMXgdIi
nNl6B8Qa0CeiJpizp8X14XjbXAV+Dl7kEPSPB595XIoPRLi01JSLX+Slgk2KEbna2pgw0wYeE68u
DTHcvYDPaq9Rg/lDEEQo8RhLj73BtLE2kD6H8KHW7cM+kNJI2sthNxgMfiMgqI6PYXpw/MhsnrK1
GLm8mwWIU/y424fDY8yKhzMkCLswM1/f6udDRDS+0C3uUIGwWDMKeFFlRBX7ZWwSacAH2Rys2z+D
u7gai0BRgR1WIjzwd9BUR1x4xzDsCluZf+/XRNrWUGee8WtHRv4zG7UnhZZEd8lKxcnJ5AEHnctm
4e0Cu5bNxO5my3bjomkxUOxZg3dftPowCxbBcjYYOJtdLhSuS0YNzPEYqUcLorNWBQWdsRGkwLj1
FJRxM7AlY5etVdvfUAYWmmC3BjSB4mZCIWlVPEuexD6ztwVt8oSo8um9hdwBnkoWxH7Kfe+m53f/
+DUKeHLSYEskUxGtcmSwkpogVmb/6RYEC30A2dJQm1wPGL3B6UtI1ng72wpH9PpNeaH6mfxOZrSx
KIGrPrdUtc5uo6kJjtBLaWV0Mew/xt0mSyeEwzmaJ2t5zea2k2bUZTrPw2p4EwCr/gGp2HGMt9ZG
Fm+VRwEjm/0d5CtZUgWpGnjJVGTv+iUMw/PYNMRcdFnuDbSjHr9p8OunSh4GsXnl1KyVU74GRl/m
o5DPRfJ3hIAbsf8Fs/pjRG1KutHAyN718/qf4bMj0JQBKFqix6TOdUzVOuyg0JmtdxxYTohmT6ps
R/b6YfLkBIOIjYqlYqwzyo7xwpw7RlgMVJvxH5zxUFHGb2T2Z0mvZPG6R1XBZYVRFRWVwHLIssOi
/WY2Bg45a1o/w9q047FCI+DHJdLWjC++HMOzGOw47jB+/6IwjKOO9dxwSC3vTMPBKoTQAEJQQvW4
0TReQfk2/82+VZkyKPQDg5o3V0yNMn6CX+u1EtLKjSvcRmc1QVaKEweTIwznXRJFIH1XmtNNMi8K
KxQAcpglLH9XahGUydF7TGHqXfHbySHbzTgHlV0Bl/hEaS281BzAjO95ywNfXrJsC4Ek38prgFgj
SgUK65HzxGLfkjP/qYPzQCAcX2tFuu2wvBcageuqBn/hja/Ob/yq9nE3mD73F44G4ZqibIYblzbn
V8UWY7P+/j0DvBX4tGfJJeotVfegADBAKS0bTfYeq29rdWTlHWizOgJbp0qFL3c6THyT4e5H16SQ
+9lhXaQYn/s6svnzTw0HzxPdjUBpFZyMqYPPbCYP7k8EhTyj/DrvsP5GRbSzIVlfBXTo5VZGCeda
SnyGlhTRlsN05qzBX/sWeudSvPx12RgDyPVT872uGJvnKHlNB3isfhjM1zzzMPyY3ryJe5YwaBwq
GQeHUwMm9PJa8WsRnXiBHygo50/XMj2SyBntBhkVMvrIBUQ0xOm8nfyQsWkv50WpbIBI7cA2wDxS
Gz5/FZHcqgx5L0ltFuslsk36Rmx9bD+gMKpDZFUzoJp3hHPTZelDF1dAhY0nUdY5O4UGpnwjvkuV
DBtDaJ2q7IO3iB2AJBplu9wRUf75Jrtl8qnm7lilXIAsrEQXjY2Qn81G31DOZlw+fcV7w7STIjgo
xOlP9YmG9Q55YdsCJawfZI26pGaG0htln/tzvePJgkLV7QfZ2v0EYZsrrM0uLI206taEhyHAhO9Y
MgZM6ufxF+RM71r+Ob5ZX92PRfFnNV8cfAvClpde3E/W1Sc+ItqxkvJm6hdleoSVeBSgTYg30pxj
Krw0bZe8aSroLxtYupERtTxNHKj7BwTnwR8A9cjT3aY2MR95bup5zMBBTJwtdsJMZxvHnn/v/X4N
zS2/Baq6N1DUJ51adUt3qUBE0dIDdobVbXof3H++pJZ8nUDxAxg58mZPtuMHLzObAl3uYoflwCUC
Yp6UCNUr8vzZdcBEKm5wLzQ/S+YbNT9eVRMZuX3nA2zVzoQVb0n3X5CKFc9pgncDKMUkW3qmew2x
eMQNlvViRVFwpwXOk/ZE4HrebR/GS0DO3mvrmkFBH4aUj3Mim+rfQKidlWXIMD+KdeI8ZqazZCSj
P6evyPeb79eDoFqIRxsUwgMlCY8OGRhMvFB0f8gjwVSpCHPTMa1JXerVljY3djbB8O+ymXzh5dKm
jZygT1Ho19hryk/Ph0fRJIAVdnOF5qPpBkEnkFLg+Hm8kobc8KWTk4VtpzyJiun17XxUB46UTFUG
knX8lJDwonYI453B2By74ULxC0JGqO3wKntrAzpJnREODNGBwRrhelvMn6WLuYTGmyU/MAKc/tYs
UqXNn+RiABTyLLSXILA87SI0rh/hNuAJSafGQEZd7zUy6PEs7PbqjRJ4iwOxA48ylibWsIiL7pbi
SQbAPPDH0GdnMr5TvMeZBLNsak5kGQ5Hxo5LvUvdfPaV6zKi9NANVSiSsStYWfixcnuPC+O/j7cE
k2AbQfSpCZjp9vdA8mMhFnRJeuR+3HcMs2g7x+VE4WzVT7M3em7QVV36gI1KrJUpGl+uwyf4QHyJ
16w0m4g2opFdDTmYCgf+bUBZ5o8sEw5kabhO1JhFi7mVgmDcJD7AGBI8PDl+bvnrqdxE7aHJdtkk
H2S+bO+pC73lVZ2r5S1OqFtnfHcCRzkYT99WQ3O7eVmrNI74wiPB45HWsgy3FlMV4jm4eO9aFgdg
2dmXGy+B2TYvvf9Os9A63IPV2lXqb+a2u6F/KkgGKXsTw1w5eocWVXzuUh4Q+QY12MDZc6XB0/rk
UPV/SSXlLUXu89MKmzJ5EKmH2d1cqU4+IGNAnmtThYCGZLGvJbrsKH7I3DjEex2Y7acxIVopgrkt
MaBefqnqvtMC6hIArAMTmIiPsS7rtKDJamd4cgvGec3V6FcG6BDaVj1tzHFB/WNaUZS9FYmEva3l
wNjdhLghZtEM8S4Lj3reiT6dRRptY9TDP1iEgabj5cLC0qU8hGKKcmUpz7xN2Sqhp7EvJ+AcB601
Xatep5bajbVLCrnAtizqivCwT/RKuWGgHnQR4CnE2f1RYc2FKT65J9+SPse65AlJHzqwrgeI+DuM
LAUp9BoZCyAjfyQR7nLmzeC1TvCFdniS9TRf6OEqoj9fPjK4HlFX7FmnD4GvjuU4U/BJH75gg36/
EL0EYg3oWTzNKe16tc5OSIITnxzzI2RGnA7gRg2kV8BzqNU0bbMxBOlsvZAMDTPlrj2W8m0R74wL
o+w7u5vAIEmBvdMlohjsdqTM8KLZaF8Q+hIqX8BGPlw9Da05XFjYXcPeXyxMPx9Tw2ro6RmubboA
ba93xBUULZtojvtmOFvm6vCozkwmZQ2ydYh8abm8M5fb99F8CNitdQO6I036VFS6+EzEBKLmb6IN
HWzVW4QvW6AxpjoNXUhle2Y6i9zkRI2MnkS8dL2P4eruEsrvKwXjRabPkbLP1WVj06bYKEpdYclr
TCB+uJeiLyzfOGdQSiPk9QWKpYcX/m5JqCqZxktsqhq6OcSqEkcnaSFHK3OgCDTTPQCkUqJONaec
1yjcCT2nNiw3KikRkwQ8pi4lK/w4UKdgkQ4aqPLYJa04S3erkBSpxTed/DAEVFtuNCf0qAdIOZd7
lb01Kr/AxQE1SKi8dDoKv6JpfjmEB8scT5DwZSYXF9FmAvgWk0HT/YWgvIH12kNWmhasWdT1Mj1+
0ZIuJfjKrveVLLRiMwTLVSR6Lj35nv905wJBHVWkuK8ITme6CnAGS36NIG9zwqbm++976B5W2ZlH
TiUjm3jy2pULxzJMg5fIk/BAMAYG3OnNtg05NkkyP7yerqe3If/n3QEs5jQzrj3i1Vah7eAXtl9V
plm+8fe+ZUIboj0/LXXES1EtWZvMxmpvArcpRp/UDZIJEUph3M+P/POekhlHCsAWTNb+0SYToRSt
hR01IuMDq+6aZs9Hj6LDOMF0wjQ9teQ0bt9sUYtEJxAI+dlhUkf67C8PNaX39KuBJ9YVtqlOrArN
AMVe5A7wCM6gr3zcARj5j8FMsUbpS67LpCIt1Wq+s3dl5i5T0P9bJFXsCavcve/jmY27pwkkcxvd
M5T5mVekspVatnRHrEgPCaa6UhWlWJOfUGU4eFz2ZDyquGWGCHD3fmZ7Wmu56MiJckEMZKTlsegH
4f+PJFxSarD+almKHnwRRmmBxZPK65zR5V/fvw4q1LeJzn7WOJMj70fVQjeX52BXuDHR2GzpvANn
381MgFcHqEcGUvJrZg3ypEqdCkvpvKPoDQqqtF+AU8xIwRoxQDaQNKX7Nh1926/o1Xomg5/ARCnk
hyF0rV7iITV3hVG42wGbc9FsM6cQ4cOuLWe4062eSzo6nF2AYSML3OJTAtxkJ6+ZY9uzkhtFwjER
bd4E/WXPFnQaBs8Q1oehpLM5NbW4/b/Hzr73272KSm0c/KlEJ9fB+eYmvULy+bRdYmI8NIDvVFJq
CkbqOkhJvjQOsCJoHtnMb90Q2IPUIbFKCUWDwnrbr9qwmpsU0SeK1TbqLflNE9/QUq6/ChWHUwA5
Ie3cEca1wWor5LjCSDuskobDWEBXqvbho+eZxvkx6FBe7+/ZdraKnvYzMlTzvb7/v3FHlNBw7wmA
MBJLTSciG0IehV+aZy6+EY30fpfZxBo3lbHOGocOFmuqbGNIdcTTbXhsUVP+LPG3KjtdOq0QRQl/
7CRCNlbhaoZYzGx7lu8rJheDJGu9Ye/Mv0GJz8P74+gdvylu9/v4L5ue1ATHUor65WmblENNesoL
Vr94Mgzb5TzgbZHzB6Wmflxl2aieoGZ2hWpVbz41zE/ykh3BajuSV0f4Jla15d98ele+ttuRkyYA
Xsp/+CORZJQ7xpXz1bIxyg5eCi7LSyfM7d9Ti8O8Ptvyna35bZSbC2V5qhxuJnVd6rCxGI5OSyKU
zVtRvS7GQbbZMPsvF7jjGqU3+EGvT5xkA+Z6tWOw1TWnE8Z2F3pAAJ9QSAcuRfHRh6TcuhTcrPke
TUB+uY6fGkGr2Bbq7dStE/9mA7CPf99OIJhuTFPSwFfCRBtrKkTGlo6DZ3a3Pl8yXbsbSRcvXDjK
pep0zlTzKOIlVSbdNVN+US8rTJK8u5P7gmAQCvwZEXGKCwm8PDmO/ZMOsjFZnf0LY2JGufuCRBq8
98OJ85PTsXb+yP9FtW9E8timKrMa11gidyrjkisdcxv91fXFXpu9dmsBvq1kZFQoTZMfLgqZkTXu
wGMkVmvael7OJy43TE5yD9FnP1VAa09PJEQ5+OeZpsODb2AlSxfXAzJJ0DI1WcULBHNN8W1B7pg/
FAs9GULiJ45KMTmEzwAjyauGR8sY48kTU3EIQlNMmVPY4pq+ABKogCUtjHyXOGjTa38xfr3TMnSb
ryy6DMkfdMCMEAHCR+FwYyDEh8jtOQMPaoC8k+KoAN54q6DGHEoQq3+o9/F0YdlDfSx2dzbh/K0h
UeArUafshEO4oEQJci6HF4rws9RZc8Ed8ami8q04RrK9vpdoK27nk+G3MvLUwHY3qjil2adi81lO
4JC6W7pi9LVVSfmeSNTp7oY2BgO1qowUeI1D8a2X33OjWThmdskxKg15NwdpgUnG3XPwSJbMuTcn
CPISh5DmRPqiEmRusjmpS89gspV2lEmnZ5ETKShI+ZfKuaF6A8c7GffvhcfOODheE6dQpibfbf55
vvFhuwW1ADnd0xd7Ym7PJAwGl6mKQRT9EIyiIc+qX49fLCqKIqGEDpfIzOcA0xHvJ74/tJJMFHq3
jFD899o/y1XluFaLoN1ZwNiZkHsu0EeX3D/ITHMpsTrnGZAZUyUoU39l7qz+OKPE/Jbms6xumPWD
9Nc3BPyATyWhnFafge0bFQl/7+3HaFaUxg0yD/Ze/rn4uk/SZeMjS6XBHGA4N6G5qVWUkXVzr/7/
OpC/iDkYdH2qzfbAoWJLpBN5GiyRytC9pCa8PX7r6A37ugl1Ho1mdFY4ehanvVSjDQ/9vFVteLIA
FUM/RR/2vpqCQst4WFKYMYISAJxeyY66eLku+eKAwH3DnYVh7WUrqcvqxNYMcM3JLKkyTgNja4h7
MCer6HF5H+i9P7wxSN8v3fegGf+xW6m8X/wp7uwgtUrcWgCQOsmuxSEMlfmAeNo/7T1wHgjIDq2T
/PHgozjgrOcsOJ0rQyot763HB0GveboATcG5F4FrGbUU35vMekaWlgfELAYL+pzQ6Su+fAAnSAlb
ELvzxUh5odZrSiytfDg8ZISCgqFXlPtwT5pgqx6RPF+ZXSOAyk9hMXNeWGG3kbWq+GoyT/zWWPyp
LIyrjm2kEBO+6XpXkoXrN4Lr/6u0IthR12p+JvnnXPR3XdBWtUv8YylLXk+TMme0s6FiMNbAeNAo
3h4Q3e9yuphlgubsihy1N8jseYwSm787H1ickHD1X6CRQW9gk5y1NJU10R7s62s0jTo7Wvy9NOwh
5xfM/69KLHVxgprB6/yO/28pDoX8r8unCKVktXybDD41hnfQrRivK4TzAn45/7iv6DeXqxzBzt6J
8hTNfIljCSExN/FmjB/KoQmxkz9EAefq4Bm/7SY6WioaFfT/bkMxKbcBs/HYmF4gfze1XAtzU3he
PNI3o4DRpvTS1xLjDKVkvq4daJgmEOp1Pu2n1cfGSae2Dh6Yc6W8TlxOqnkBOLWxrg4QGkY2C6lZ
TD89sU5Wh2g8MeFSZX9mjYzD9wGg2ni9RalsJFYJP+QwNDO7JEVlvAWCPJ/2exsjG2/RBuAsdrOp
hOpr8P3XA1qlXqT3uATFLJXe7sMkZ9/b2QrCbPGWpmihKIKPuJkalKxb/tFakmZrfLVkZKFpH2A2
qgJ+/EOzlv9KKzXtYEroK0gSxgcWR4CZuQzOLxdtOS4vptz2RyeGubCjbHgQ2ZFNG8Lre/XQa7F7
1KHs8VYG9cDWJKNz3xZuxDUXRpLiOT4/6g4V46ZOdVrQwNOk7NN8TrJqo1FOBtoi1ZZTqgDvWa3J
tc9kkxK5g9JyolkbdpP0l5g3yEaty65TrAF9DL59LMrWOMaYarRt2+8jOtX53mCpR8bJOm+RH6ka
DMlEflcgy6SpR7tAB0j7b9XZ6qlU7Qd6ZxTlyWdKDgUVD0qXo6IL2nc4f3eaUihotTO6U8gCLjGk
8OffsT0DLJq9cCWaUaIeqwEsHXpSBnJBmO3HRz74Um6Q4cAHNrNd07YSFhNrqKCFxddyR6MBFt/x
jsloCSFtH09/TsoxNM+0j1wEUH8eXfK9zxj2IE2WQedzZfnR4CxJplsZctSO+K/VCr6xmKlEXa7j
kjxdleYofQ/RpWPYVaeJZLWfDINHdkWyNC7mFFaSQMkzZLW/QDOZBzPsci3GR37CnMpUixeVNxQo
mvHzIxti1f5fz/xLL/bkCxxgeUBgDJYn+lHEMEEFSb1aSoTkG+0pECgBqVAWHNyIMVsdBVlhIaVL
jxs8A5k9bFZARrKwXooCXKEwaZ2rxLsFvGqDjbHKkzCglvDFQAjXSpn0hikOSxjoLwT12ATqoDCA
3oPnO2ax7h/+MaTM1mGry6GVvTO7feQwluElbq42r7P4s96Ywvp+KJssZ7K0xKSHUOBxvkLZjBkS
0PwH1BocS/FB4PUUug/vS/9ffBZy+PTSIZ5xq3v1RTMDLrZqJZ1b2rlfumdttR/zvCQSeT6aQPm9
i29VLih7zy2SC60Tof2K4o5Olpd5t8jTCWNUYuFio339eJMU0ajNvEhB8R4fWIN1zu7Stt7sqFBZ
pAWktk9ZGqVF2bYxMOjHBi+FHTIsN5fuSCYKmWe4qX4tpUCkzjABDlEX1NAy6Dexorr6LmhfkEBy
A6vWPbKfst3w6br288j9ikORdUF8Oje8UeAGiThVm7YL5PZZCPF6/NvmZX9bSlRupdgCX2d/f8NU
GNe1gl0rdws0NGKcP0wknov3uB5SEY4sed6b7wOv8tlZTWzFXYCz5JNGtp7yFC5Fxx6KcL9mCQoi
4L3Yi8FhQDyXAiotm88+bQOy8+Npt0VheneRf8EDAd5quzQL7hAUPApqrweoL9GJ6GsvNF9yvim3
g6ZOT4vmePy06RTlPXb/Jlgnqe237x3nOMzrO9YYi6InYQLl45GszvgfScGTE2J/QpHB7nvnZp0j
Sfv5Cl9fk0ltOtxGBHyh7k2C75mynk4mTvhGmvzL9N18ulqLxjpk2eBSYFP8arGT9FTUQkdTZbQ2
1XkdK5dd9s9WOIfQ/ud4WY8Qb04S77FOjWJ+nHCPp/tMefV4hZa2E5wwNo2pHgeXHEJ5DHQp0jAD
RyC4tajTtDFCPnh3KHL6GfwzQ3J2ONLiZDdicTZSp+gLs86DbgQn79WaREueGBozCFHPLCDRIjKE
iR/W10mgv1RCSr98hb0jJ/CHLycaWaLL2FsArqGKJp0tFchq41TFuGnFmTfAYw/v+SiPLpW3UlXu
pgYQSCIwLDuzEMtvmKkk/ClbeG+je8g7WbARiiYTea2Ygbg4V7xEXG3+qzT0U5+5n5+0IvfWtfrt
jEiliiynU36/Y5gFXCRDq/FdQNIwzoY2eXUULYPDieqV9Ri+8O/xEpYgBKlTdN6NL+zaHiO/0LP/
J4N68kZmpRhRI9d5GFEw6WBr0IZbsBeLCf3L1ETXpUApnKIexUAr72DkKs8eSZRLYrg5OrkDusN9
e/D4tU65/DY9GjREZI+brdl5dmwmgBIwcS6UCvRTwx2tzXS8lefVoOG5cK1kuLO6kW6/QO9c4VRc
NJW5jee8pQcBASbjegHra/lqltZIAV6LaVFDp2e0lJfnzIs7uCsrsnZh2QJxjg11rcqllDRTE19X
6LryKn13/PUr7WuP8bOx9axDEZr7KqtEF5JYkSuSm04m1chnMG+aDFwg89GGOaUL9K+6k7B2tZJP
r+h+13mD24R0dzLCebdeK5o5ULuSKk/Ka4/oNZ6lAbo9CWiPDi9eLGzkB0p707SbLhWVeG2LCvd3
oya0PgVSLpe6epuJWLHDMLpaWSgUG0c3QuxYa9ukry2GaBby5K47+R+P/9Vi9uq0qSIyW+B+XPfq
9tnuTKh8SpAPutI4pFKDmEWkiP8OgVMs01GOJfi1D1iNeUa7gFp/xJa+aA8dCuasOHRU0Ud4uHcS
Q1KD6B0AYZ3PSwFUo+DegmQlNM3imoBg5S8K07JXnjT1y5EfUCZMMJaHiVnd+MjHYi4WB7ES14P2
EdXlw4H8QJsorwP8tjL91+mwrCKkg0gw4mLzzle80g+pi8KzJMkYf0ALJDw9QxAMpBQbHGxw0IBp
RgAi+zpeTIivPDMPBAbRiNWF5c1yv7ECk5xk35XbI9EgeOTQAvIMJqXRHWwgme69/eejv9y03foc
0C06uxnfqyf6kKXWnLgk+AX9dXOwRc0CftbNN232/DwtW+hhA2Iu8Kmgn3xur6D4dx5r+p6H+00o
ofi6YDFvHu8VIje96LvgdLs75489E6lUZqek0+yGR1qihloY+KNgYvsDR6REs3332gdBljLSJPQ4
5Jl1nK56tV3awfqz7c4H9p38Nsqbalpm9uFf7ghHJzxaJBnWzfOQwXukJZjuMAwVHjqZx6KkAkXy
kp9Zx+nXLGW/hdJRTYiYNbo1SXnUgrlPT/Whl5KnOqFeITcFIet7L8YxlCweqc4makbLlp236rkM
IKkAWfx2ImpBc/SFtqXv58FzY9XSYgTMnnXi44b7KER574j4hjnIP32rSeWYCqTLD3bnzrO0Ar9r
bzBKxo3V3+ZLkgJTWlSyu8nH8SWPQPbwf1sxITuA6jkPsIB30Yx3lMso9FlR9dYaDMMROwaxAUCl
Sy+dlh/4wmgVfJYHazbuzxyE3oLkAuafTRqK6dae5v1N4AxOuEdq2Zuy/J7+AZ/GdmeThyFWIze0
9YNK+iwROIeCHV6zVr/LmTCDqQ4ukhDWKOTCt+YeqJYiNiRO+zQ/Im9Nb9ApV7+oI12upTMK2PRA
E920kyi4rsQFqvgeSMuuVjHKQXeX6YlpPb9Ue+4dK/M/4JKf4pibdue6imLYDKrX6zMto8JXqPL6
fzcbn4Zk5Gq4Gk0eL3aWIFIt64UGgssfoXXAVXVB5RmzYWnnwdRhlWn4l8Izr6v3R8JHQ8CMYqvQ
A5/0b2LwWGsB2divVkuQYDR0/NKOxfLqDZuM1szlKx+EAOpOf0mVU69M3dxrdoTeQ4ltBqYGrIm6
4Pp0hcWI0xZ5hd0ywL4V+12jQMb02pcxeFpvuOoiwWZ/8srJppa0KvIAUisgiyXQ3+g7AKUMcGE2
p8WKhxQ+VYabsURiJm5ZmTX2WcOedB2ozR1Epj1t62vZ8hVtjCfG6J9V5EqlLgTQTB2GUmJKX7uL
imaZPtRJxw2otAQsgsoZsZxhi+t8kUOs2jU15GQmWvy+Ya7TzaQSKsw+gjN5yruFMi10i3QNE5Tn
j7JnzM9KmYXVE2aVUHqaX83R7WMutcgJyDUAbjpB0YCW+5Op7n0/0yTqzsjkpkbpWG0RXaTpRj8V
lxW5TwKSlAP3afnM4/SOmOXxpmm28CQ8DkB+qGrEUDx0j3cuuA3ZRF5FXhxKE2QOdOQx3/+XTPp5
yvbOiXcGjDOjvxCqaurg5OCM1xCPhLsxomWljtlXCAvK1GsSu0188i7SwRWjIe0x+eOZr4S0QJlY
y1NxnLQ2+azGOyDYQ3qHb2tzolVECbTeClCsGIZJc3ID3H5CQNOmO4VHtzWzsDippVl59K/RAbom
TWOseWBNP/0ZxoONdIeGFN4wgN1qCXODuHW3pZPLAP3t7jifrXXmw8oelezsOGYFybrjUacUOON/
13RiTR46LhoQBNV5D6o1uRymu64z2Liyn1MFJ6Ce8MC4XLk54igsGOKnK0S8GhASqdqEslcLwgv/
oHgsld/e+TFiT0U4gAxZnD1qAg5glvRvTTUtIoXtiCQwxvkLo1lhulepiO/J4xTRasNccWgZx/IU
v0Wr48AXbR+Sd9o+QycTpSikBLsCEceg740+th7A8WDoZV9IVyIJEpZa5l3uw4YaI/Z1cXwH01B0
OywvUkxNF5MidjYlNz1F3Pr7eXA8p/Wo/6P/Gzr7HUa+No050MRoaUw776ScRwKbu5vZmYoDle+G
kfgIUDg1RW9MLjiupIGjuCYixeDSXmgx9quBw8I9qqAXV/L5uWY3TNspGy5MeuZLiym0YDVgTBBY
gBC+xs6eR367vwD6indymhVFsvp/ulElqkW/1CyqqxXkn/UASeTU/MZdjespOLM7a6bOSmGPsjEn
tYlozU7NbHS0Yn5v2GJ4DKn/ECh1hSgFdUrL000h8sDQVXsY38WvPRvuxaB6gW4nn1hmfwsWoNly
HBg+5rFMI/fCalhG31Le3dnBu+xWnW32Ju274hT5zFtu+VQl5VvCB4TPqBz5WL55fz6xVw3UpFVL
CvDdAB4hpOnn+okfYDqDOA4Umtja4BPbw9OcevUsKMYgK4tj0yHPkmB7ruPSK0KUyh3wSQa/JHWx
EUOO1El5neGCUSfbgFRb3fZfC2Q9+/paDT+nDphOUP3PdrbqKMyrpAXjm3Ox7ZtxXaEQg2pelMlp
86J3EK/Z0+nnsV0uotWhaviGXM/doVOW0b2Izqkw/s4cuRaOcRUSNo65AK+stx5ab1MU2V5cVoyo
U/koV4kW3AWMTEiUgeGuGmr9sMf5CZXmoOZZvuV4Clal6JLFWX8wRbQJCWW1LGrgYj1E/PAGSQGb
cu0BYI/THf4ezv4cmmgMRNytRn1nDnu3LpQPCXANxFdRxPN08CrVoLDD6hBWF1u4UiLlwhf2M7u8
HWAMD8Sngnb2RmruSSWIwEx76OaY3UkG0NzNIkumdZWtcoLdq3snXYGayqaQ6AaSaAivvUGCF0It
OxEYqIXJv+Ao3fzPD/ohQ0ulB3orJzmq/QsiPCVVAvJS9C/4hUzpzV1Y8/3X9x4E+qm8wg6Da7Ew
noxiDy4dkP55t5LWogTSun+TX2gJmzkRmxHROQbjHTLj0Lfn8GW7AWUDrhoLp6qt+EDJ+/Rp8+Mz
er59mxZzJDt/Wry0+uBIJfgo5fvMYmT8nXOJ6oc+zS5uhDFqMTbKOrMQrJ5RuvNHrew5S68kwN1p
BQLcAOEcK3uRf2ZJ1QLM+uxdq45QvR+SSaEPghnaz8mhAkUIOlbr3eUqzj89E+4CajH4Ba5969CL
79mCbYgAX6pgs7LHUb7gYUC6rrdr4eouYg2n3T5MEDP9NRBqqXvCMyfvPsxQ9M1wqXf6qI8zYMA/
w1v9tljFlVuLNBnKSnB/YueFYWiLFuhKyModL6DLIVI0MQdupCPSaXuHPo/99H+4/IK02rKyFQz1
UvzQ3Ry9XJbvq/1s6DN8pNhxmIeJ8SaT3QF2smI/QrT9t+Dwc1q1EGlWtYD2qWoqLt8pgLMKLnua
PQWNv9LpGIJuXxIyDQEGDeklcfrA+ZLvWxq6FmA+ReJ/LgNlqUl+PJbw1iI70GSVFcsDpwUP3dp5
zMvmN13v0qVYD1e4HzspMMMGfECwiWRl7bYdJGvYIACYdXyeuHG7/fzP6G8v4b8Y5RL6gLLjnQ9W
MzpvDO7YLVkOCqgAG2Ue0rNNuv8bg8nMGSixQKhjf/aasM0FGE+4bB1gNtidIRQ2HENb7/FcBzE4
MBS9gQrrzs4sk26vwCFe+PVxxTyPaavsI6C7bb5K3jgxUAnjflH59y6ZIDMpGjP4fLhC2j0Qw1Tc
5WfSg/5XdDhG0GT7qLKqqwldICgiRhdD0U6aNX67KGspFdN6nDLnyq52Eg5W3WWgMp0cWxQt2N7j
bXH1uPWUuyvH7rJfvs1bakjHVpg/mYGcPm4Upvp7nLMK9tZyqsY4kgbuS5xv5Ttd+loWtv5Uyj+l
AdiqylorxudL5bbbn8XX5gUYH3DapjEdj/rCK4U9ASkKVcCv4a8cP5beyNieDB8rJxHeD9ugyK1J
w2UtrrUL5lxcFeg+eP99Ck04P8Pn4rRnCHnEhDQqsq0ddH6qOgV2fv6Mslt38WussLV6TTyH4+er
0UvykHggls4GG3rqVVGFLSF9K3ZsPIXiRM3l6XjvetGfC5pmZJgYaRV92CX5N4ZrXXgpdTq58Phy
oYN1P/xi7s9GwGctaXIH3QghgsB1iLuVh9rnp2Yt8KSDA7JjOAAVRSopme9WNiZjlq5p9oOt/ZjJ
vNzVzAkULvW9zMzTwb3DPTpRaaYD+DNQKkD3MICyCQSqzHCy6UOtnVAkHSphnA1TAdbBVoBKIp3v
16pERDmm8nbJ7zaQoxnDc8MK0KxGX959tNyL8poXEw7lu48uo/UFpFL+SMzhXi537/XjC4obSF5u
WPzCUTk9e/dXYQ4o78+un/dCdZdWEcFOmswaWZz8aRzb190ltS5/R0sagzjnBYrYweY7dmXqCoAT
xVBdeHigTwXLVRNDs9rM9npfT0Wbo1+I79MSwCXfQe5EI5GP+x1d9Y/enbgJqTkWF98ZLgzfwHxZ
mIdL1S4beqD+k1jIi2H9yhXYhEiB7V3xFfYRe26DVNJ0sh9bSSWZvvtFiV7tM8boQtG+oFf+23am
Obb2rZa+Ytq6hYawELg3Kns8zcXk06Ki2dPGWxtpE7o1rlKWT5xC38B8IvkzbvwAS8azZHUIOe8b
81//fxAKsuPS5kWhgO27fpGOBJ8TwIImZrPoP1n2HUhx42u4C8eCIKky5dTGr5bmW/MmjGg0dZnp
XkbCNAxwmJKRUv3b2mkq4BxLhnaRuqLB7//c5b4EuJa8HthF3Qm/ZVdULlfnPyNnvcUrlBjNelRF
e7guFcoZor+EnTU4i1AivMNTswKHs24p1JPODlgyqhJDjOJppR0qIEHvYbk24eidqEwlus8qIwqZ
jN+wt8u9GkGQ5+gdIvwtJl54kqJ4UonP2kQN/eaNNRAS3x70Gl/SK3J9Bc0r/FKOROCMOzhj6WtL
M6CCAhPr+Ey5ylb6kyCisR1OoMChe+e8GwrOY8s9Oq4ehqocEKdjO1oXl3x/T6/yu39x8GpIii6o
CHpQ/IWbaNEQG/7baHfQ0NYSQ7dEXk2Hket16wHE8WCaxjsPnlhdwUJHnA5ZQwKwj51K25ukun2a
dmkmTav6FF9Ytf/hkwQQqXBgkBoMGzD4MwwpHe1CWtaD1Rt1E/OECrpmbPnO77qeoR+d3otUI1Ol
SyQcCZC60UveSai9/GhcI5P7ue1eWkaIFBL0IByqD0gtCCWpLtqgTmFfeYSzad0yEuiqzgWfa17m
4AcpKacJlXtZK6yqGV3dXY4P25VaOORmkt/u8G4ibVklXG2qWeObGZMauYkt3fiSzZJgR+begwN7
WCDXKev8djZtq0+WH6MawRKPqbJHNvhGquVFgBUXg93aeQzkorLJwE9cS754nzErkYmBzQiizT3P
XXbEj//xM+AZONCkTDlV7zEuptovPk34rbh/iIHcK05f13XTN9wSgCR5j1HdpcFHya20DC+WDNfj
0ISwXeO118d4/IvSpNuZzXLCkSeH/gifYI2WBdB04RvKB2HRGVs7RU2gnPdERzUhc8EVwZAKNFD3
uQEm0FNjYqB4L63R3MYJkwvR+8FUPCBDMX5ixCv1thnDoFw3+YspTkqN+7AzeKJIKI9fU8O0yYhn
fZ4hBxpuP83W6QTd1b7lmwPVN1ioftPuqGJONhC0VUAB1NbwNOyO0kOfUUguXxa577SGTJJtvgaH
zq8ZDr2OD+Sx8Iu9bhato6+KxskHZTHVm/VJbWYn1sUhRyRyskrsLarUuhBYnedi8BDSlCtgck8/
nxpy+q0Owa67Qd4QdZ2pGYVbvQibeaxsiJjP7yIsS+Qno/S1hTEf/YTIeO89x7A1sOI5NlXDW10k
wdVte+Cv7cibMRRUZOIaXJZBWh+UfONYIhZ1LZFe3c+IK/SjFQCWgJZrHAKb96neHeST8sFn2RUB
GoxqjQS7bI9li5jS6rmWjG+UaSXvpVW5mVAt1B5feLub9v2yL+Q0/8wDRbHKCR5we0DH9kxrQAZC
LTUT7jK4w9C23ScZ4JlWIB7JL57cuyZhq2Si3H6DQm08CCUfX3fPwa8RDCwLoUlv/zc9zYg7MIhb
Jra5LfPcMv0YMCb7veD/D5NXI35Nz06OLQ0bFur9I/p02QyxAm2bkqqY7Ey0aMK22VhMifp1P+00
lFrLbYdUwvd4B0QWh50aeiCHBNmbIkqZPqTznN2GVn8lG3fwklb1HarKPyBsg1antDMTfecDqxGf
4jNPAt0mH18QEYNmfjs4HN+ni48r5AgfzJkfflYrIVNVYtY2EHcEeP90MBN4aiO7gIPUXVnNlsIl
GAyMpT33vpz/oRHJrb/oQeDRmVPmK5tdL5QwOOAYEPZwEqjabaE+hnowhhxO3rpOVgsbH69OV6tA
9a7DQK57ZC0/lLsTDdnjPSuMSWAANpjo4I2jgwX9hoIII1Uj9GIPxtVnhq1wz/H6q7p/0cFGlIDI
rfGBVuSEKyoRpZld+RemtTJgfVrOd8nflhr03hH3TsrjsT7oEv9Z1QzN8FSanLqCFHlUpUydUD3G
WgL6dQN698jo5qPGhSyqKfj6IAWPoWi2F+kWCk9qJZ7xLjWVrlbWaFb5BfvtWDOR0Vy8Cl7NK+XS
eEEHG88V5zc3AQFuwerckuA6XbSIqdBjZY92UZgtiFovEKYIGzI0ExrS6XgmTT8O4p5C9zua/ZCT
5MsXZ22oyT/sn3Jiqt07Q9B2sz9tJJNgJW8GOGqGBjeFJ+lMlxjEB22hVEiArMp3YGWpLj1aPfy4
EDNVJLbxo5Mvxu/zJJl9Yhf05t6dOziVRL6FCa0ScA9X35mH0qI5l4QwQbTuOOj6x7zRzdLHfIVs
pAhUlHGiJ0qI2Hc2CN+uTaoOLAdMDNABRow+1CuVWuj+YHZYeXs67YnrQCkLMWQ0XSoJqmi/ZXcM
Hhf9sBdV07O57UMU2FchsA85uWSYq5Zy6D9ikwBEaKc5UamINW+px2bAdQUcEYZdpDUxTS6ySn17
0TBDE/BrtwCucIeLQtLITE+mrl6dRxjKtb99MCtvU0wNkg8d361dGcN4+J7RhaV+efgK871aVrwJ
VUU/h+GD0b6X4nzRsZljR39S9aR1XNLP6Ko18GGsU5ze//ctGOVp1+TNiqrdrbNbTbhKayZW882a
xx9la+pmBi6Vw+Kjh6nv8h0OOf7KwJ5EGMizX3NzmsUqU7XJiGG8BLC2DLxW8Mlt9xCjs2i6VWl7
wtEvozTtJBIT3uVPdhsgD9buwd/9F5KGZgSD3p0T+GVXqOrQGH7obTyM15hZ0uGDo7Ee6GtCHUOT
+V02wIwTR0yWMBikRIFEteZF6i0PL7bU+zdqPf9CuslId7YrY7k40dJ1BCUlqD+hXcoboYBdW1Yf
/mhHRNlirtdxRjFlIOM8Qy84bEIry1o7vZiDgfwE7GPzhYCb2Vxx+X1PuaCFkh7mFPhO4FYQLxCM
MpzKluQqMqggw1IEPSaSZDqnexUS63gGNt2IS+f1WaK4V9ynR5newx0NE/rAx3+le4+yv8YWwmPA
xTXMCYqzIxKHY+GkMvPciJfeRXGujK+zZNkHHwuWhIpHDlR7iD9+fabuiFahYwZLml3TAQJ0eAp0
saDKZKnXMQqihKnOPzkz9IRPj2btFKciEDbY4gglwAPvgrXRM9DE+J4e1dmaxzmxARi2QauBIErU
2x9RmpL6Yv3m7wedKGqfBebK2j/CYtLVukuGDaGvmMmaIc1hF/OB12AQZNjD+jTfEzQmrKNoinFF
BqTdMv4XOvu6x49u3T8wzHm/jMcx5lRMYI+FSeo9G65WVzdOtQVhUR2TZl7IiN1uSXjPGwfkiY5h
pgghBM5nZwarxwRH9ykXVm4TEd38fOBdZlgnRg0rHeFUaZ7q9edlYA7u6EqRszdL+cis9rLsgLpE
sWtgFupJcdAO03jyZOC9U1WXkGBI1tCwnUwu7I8gB2tKPLGTcIbcSRh1AEOhx8l1s49dLXJoN6dg
WnTW3BZ1Wnzx0idyGvMfFxPD7UngxXEpOJcF+KQfxmY27kfbbWfyyaXFsPRjl2kKkdE6po5xH7y5
hD127nSqtp8HcIbYpUQ/LMWttVjOHSRC5Rx0jmf7THYANA4sRvqpa+6AVNRYn6QDBY5zi+hNnaE4
1x2sU7j0WYPIILa8wufP8QWHRl0jvWOoBM7d2zLgGQcAcV7WCYMhGFliMNIrgC3nix714ItB4SwH
NTb6npYJ2yAy/I91ZXwewxkqXX0d2hcelNL+MDOhokrLI00dAFt3FjDo5W2XKCJ4OqVnkj6a9hPz
T1JBnlv7gd1/y7VU/ziX68TazKo5CBRbfZwgFo6vbHUNN6OK+no93DIuT8tpW+GwpNbfl2PSrZ8s
iQQpfIS5skgypoHWqJ4AVhEZHkTl0DOhuEBKjVO4TI4TbOxkhyTVBnPvtpGz1iTaL5fStE9X8fTx
q+1FLjL/iuVSl0DK7jy5m6ArcJvWl0SK3/N4pfw1oTIkyY6KF9lzbzDOk0EPx1J11NmahZi9wdpM
WmGLh+b1CMJ3Cr6yj+0wsbf58jSfizmiXaJBvQArKEz6/ruJDrTZqQ+kZE/ulyRrY3+GkdbY8vWs
EAlRt0AxPiWzUeoxxmRUHgf13BTPoOOytA5WsV9o98XyrcBc29ksafgJgPkvUOwcu9CgxTg4qblR
uBi9PYjk86JwKIs5Fe+taTLl+FAePR0bWcGMnkbFVGkCopIEMJtDfQl374V+p4Zhk51A4gOXBpvX
CdXJ/Z3rsoPWC0AHJnmuz4mivq/gfIZwQEhdzqaXJsWHAFiwqRhYuS807Z/M953jICm7l4po0Hp1
necR9erbJcMk5qwy+nZOr1j98u+82T67b2DR47+SLauOYLQPFkCWfUS8JnqWxSOhwxF+5ydHGCUB
5NAHTMnzCWkRxKewJcxPhKc83zUPH7qII5nb3ePEKQJOV8lK/UKcV+67p6Sne0jMB3EABLfi2URj
eEJJutnStpK4NyWengBspTorEu3GSmlX7vBpz6aIxB0Wc0JHBhWP7tUgPqOZWwLW5pssEjhmT2MI
V6FnllTdXLSISX3cg8F2MSAMvQpZhel0pcKIaMj70Tq+X69YsIegTGjUO3l9yBcOjWU1ZGz/DbL8
ooCSjPA8JPZCqZeU1PSwcdTUG7dqStJbrQKh+bQKSBPizRh/7kX5qfIYVolN28z4B1rVVMQY6Bhk
iFT/vajLlDjae9HFk7mLunGCIQsav77q9KAenv0YtOeXMtjdShykEaF73BOkwl3ibarFsSnr+dv2
yk1OOeIN8re57pjqQJdl5sd+8ZCp2TRKm+ZR089jbhDXJG6SjFB8Wetot1Q5Rop8StahFfGZdcV8
ndj9WJ+4vIoAPlfPVk7Xou3mBr3YqXw9FTTb9vtUkc2iQYyHJ61xenvOeytwEc6Sd6iDyvsf0cWp
ECXuR5Q6Hy9B/RdZ54VZDyJ2ZnPeW2SUl4Kdj2c8ibokfAKyibzJk0iHiHWuxjYlQZ2cYaHGYFY1
ND4Y66TAh1qez/UtISB3UQzkX57i98KboVP27etmXAbayFpQKX1LQXOgJv6ttnzLgx1qdEay76PB
jzIdQjwBy+1rzacOPhiEk8Lxy7JfspiLC3o/uL6rwN2CIz8zxrm0be8AXNnXgAPaJuhUSKfZLpGf
iZ2OeMouOGDy4I3bz8sLWKmgz6QqYWOFtx7ui4i+herCQrbqEHYYF7ZKEhqSzXaXkNm8CTuO3ia7
pmGbxmunmTxEVFoF8gj1MrZlmqM5t6iqdA8eGlOGj8/9G/9fv+v+gi+7OxRPxtg6nAxhAh8W6vws
UKqcnFWgqSh3DJntvMYGWZn3KA2jQQH4JSwj9iKSXwR8IilnzASalbeQeBXCNUvc/8oFfg+n95se
ZoupWWKsigfeWUPzRlPQ8lV2urZdPCQBLk0LpqA9nF2o/bbCCD/8TZDzzqa7gdJVPyATpPP9dY6r
3VTw2cSdDMioul76MGL94Kx0Aig/yuMMMpxOukIuP0sIL+9OfrsuOuk710DEKyvJBWVaj7NDYWn6
xh+Oqb8wDtRpsoV08DG10aE2/Oq0X+lAwCMM3a0H3dGQDtBJIYxC9Zkmtve75hvAa7+Hk7+OGr0u
HTwpcBXvWMf4l90DzzVQxIyDwJ6w/7lNXZjqIOwfYk9hGCM4sfc6antiBomDCDDUyJb1GLtqAbVv
15D9Zfw9DR1OzSQga+VXPzg7WIRYrrPNhPOcRsMKJBY4YATCGkHwEuQ4uDM3SuN2yrohylFitLU9
Yowzn3CFiekMXJRy3YWsvVoSFjf/Zuse5v1DKaVab4OLXHqVKYpowGY9f4XFYRzWdi+MMq4inDEc
00HzHTLma0G9E+wpcX69NhPYkKBvVGpOesDwW+xTyJqEZIozX9KXXlz0idkKta4daR6KvxeLDqDT
fkpPtME93SGlZMah0Ci6ZbkIvebOYo8MVdgB0QEKYFSYFMpRjjHGK8T/68wfKL2iImeWUgQEn3D4
QhZ5PSQIuaSNxbO/H6aKOh3Z4QYSnzrCekjuh4AH/TDQB8QEbuZzFhd/nSm99xLrI0atCIvXi7q9
RnhBTgnKOgJoEJKDR2vArbG4I1AYnDNQtEuK1gruK9KEQMkbH/xs+P+TIBUfTrjjKNWGRVUcTi0Z
GQQ5CamjPEVyzmFp6uossBw/0dW8jPs47jF3S/tQqlR8LSMriLTJBm6w/suYY102fElxiIImlbMZ
P+SbYC0e+2gzXUdCcc4Uvfmg3wrWO+ZOpqeuRRstpItxA+vHdGBvnEP69rt7rs+V/4TXzomoAXMi
MFdXFVl0W4QIxbF8NWXGSUHLOcVyQipYpOjDJy8GyQ6So3pGTfpnauUhNG7MWb9EiZfO2TpavjmA
H9oIGbne2klbuXdUwrAxnuDP8L2/03U5tr9/gew701Ed39LKqX6kQNW42eEUjt3fgyrujCUDDloJ
j9KHKTZ+f4V05ggh/u6ICbTG8J6TPuOqAjKU47Oz65A3ieLZaocX+sUFIVSM+rz+kNjNZEsaUO+m
8c6rJu2d0KW/QwRgHQB5W5a4aNNvUPEsV8ZN9+p1uQEteeFunB0vpx9Voavvr+HCQWIJAehHeI5q
WUFLS5gnYQoXABFaevA2fEDjYdwgqw/yZ/M7L4qrZ2nrfSDKdE1CaiJXguN+fXVgyVQxOiNCRee5
L1linDlu2VTPFiuJlAnZZevNMNoFVmuBAo1nsgMZJkCFDWOIAqfqSdJhAk4VIEYlSRJFbujTJyKM
zj/Lbf+d7q7JHq4jQIZtZREkmDBQ4o1d5xBXzlHbruS2R1nYg3x0QypgW3ez4qlZtXZK1QKtG0uJ
Y/ztkCVtWgNhXFIezcvEv9e+RM19pokH28hBdgfZlUyBtU/wNUhBuqD/aAClR1VFfLS3fLcsa5w8
mf9ILj6jcvG6FNUc9EFSLB30xBgZ8ydKvpvvVtLJzgOhocZ06GtYU+geSBnxlY0glm9f2Uf9V5ZJ
w0D5YnzWELbjGj4I8gFI5CNDBiUFsBrLf9vEg40O0vQXWKLaA0wQcmNnwR45xf5DnnQPNI4bR5DM
5YRlIEjmTLy5TCVfe6yRZFkaSDpPC6qQOzraulCAvv7Btqk1C5mlbzVLIwoEQ2Ah0tjQd2GZgtJn
gNaHvjcrmcO16hlMsGA8aUXaZ2Nht09kp9ADjs3oBqcpcvCvQmnK/RjeOPLviQrEF27rJFPPA6uW
+4v0aqmnfi8KxOYMWVbCgL4kQrmGUgEmHbTpafTC4sPL6WxgBB2pDc1uU+lWBUlnEPjnzdY/A3ML
JWafx94m94qWhWqcePdC9SalmF5o8KEFBLycLHc3XubXaH187Hp/oTEzPPCZREEUzZOYMb1VuzK/
7/X5ZX3KDGD/6R07wXcCTGQHAz+PMnHtgdZny63kRhoKcBtLalf4rwt1V3vc7ixQ+bUFRZJPONug
PZJI4fnHsxjUQKtFkqlsJbShVgxZWnSX5hJt+eiHU09mws5rPIUyCiD0He2ox/q2l9Dqh5w8VfSY
KLsMijbhGOTLFqMFD93j4JDiNGizdVB9uJxMncmkXB9BndI/+nrioGvlFT/DHcFcfaPZxgrCHZPU
7OKbjl/jrSmpAg1f+lG/FWr+bV/a+wrh/LmoWBfhymg4qst8mx6acvONGMXpwvHu7NuxoWTqBd4Q
TV1fLoIBhi1ImfAF9Vx01/LpxKPbEhq2KhQjG48/Oz8xCPi5X6ZMKW/YRJHPtM9rc76gK3iGMaDq
LMlih04uBPmE6v4sXsllk1AWE9xYenl0QptRj6kf5hibJgYycQCaDhkS1d6lIYN7JR1aMcMgFBUd
RXEFfx7chOROTYcHqT1nDorJUast2K93hHCnYC6/8fSCOHk+OHb9Yj12+05EcWIzqVTIOWqEAQqx
4aeSy3HyS5bK/7b9oPqZkAiVnJQmqsedH2zuraN1DXFq6j5cWbUHJSDWOiIzZArPALZejPCommcJ
diRo99/gTjg4cAIZJExSTyBrMpD0XhRrYjgMhHXVp4eR7OV1ZvWk6Wp0ZSOJOMwnZglYDjUn0jif
xVbNXvBIN+mkYvPkrJFxv8N9jA7mM6GcP0EzswVUpxzl0Y/og+uQ3Y+0xBj7iocwcGWVJyQ88Ma3
h7d1q75SMYEc1GhXzss0y2zlC4nhiKd33PXgbaPNCQwZ/s/EqQaEvqSyURuWUD4Tt2Us3MDdkuWN
xp5bjYpYYoxDOzzd64Jw/QEfnXW5r3nzzqaIh8lfASlPdWDPAJ8Ger0pGIqkFUotXVNb+avgXeGS
uDZ/HNLvKnJWQ5gYSa5rEodJmUvw/gZE7I6oD9xUc2Bw6oBX1C/xF1Ujd4yyuXNfOjrsTAJGV32c
9yOqVxjfQDk2cXUGfPbcdJFP+KxzGkQLB7dnWhLMQmlKSyuD2rf8c/8p4mqhYODe5Gx9CQIqYKVR
f3AANDz7nKO7h2tnkxJh2rB7R0duFkW6RBUKTSwLZ/6KMh2qPi8xs2B6LIc+WI1vQMRasttqF7Uy
osGhXDFul1tZEAHYB9O683tBNeiWF5siP//inanN8lKmsL4snYCNpWvjUt2kzV4nsscbLSqSMkck
UOOnQ5l3vqWFiuBEeuU0nNIiLX2oqjnWTYBO53EhIhi8alCET1dEUpLUaymJ6lyxsw0pW8H11emb
hGcB8FdRw0I1BkpJ3kBtJeJPK4T5blAoiTDkInq9BXFRSJnXknAZBIhj+3tTfHVxSOt7WVoH4Bk6
j7jq0q/xk57DCfVH2S4CFBwLVzHGfWr16522hk9F0Mua4/BXko3XZHHOEtSXqZ55zEbRQmFo5PRk
blNYjIEn0iFem2xYsuGvZ2RksTMSL+2n6dD+ksKUeWLezIUYn3jHoPPs4lrnzogtraxtf6Ws9/QV
EEl6DLRzuoFcz+zwrCEEnqKnfhQK1QGwm+/ICbFFhgGR/iNK5q7UbipHvTtomigWftGMaL99LMDl
cUlS3F+WOAzguv5D6W0vxIeaJj9SJpAwJTEgKukHsgCdQRyPyvAI5tADdLkBctnD3ohdAgUPEt51
cC96b5PKBZdL6gRKeC7aSQ8gdb/Usn3vGwuw6z0bzockHFlReb9EF5O/Jrr047M9PUZVOPGuTzw0
NyKFJppovjCqRMmdEh8u+ehSE9+bBrJcomFWN5nP8Et5hcDuJILqJ3UQ8SFMhxxZWSrd5dHH278w
3tQ42r2MliP8wnpiYCQ1M3VaW3dWKwMuG9mtreQFYNLHZHUNrgpcyjISnSfdJkkyg/yeeCVQMHd/
hOtzcNka4JSel4fHA6RU1O8PkdqbhF6TeKoNL5B/30zZJXmiiIbbniF9NgXbk0qdcd0nGAYevubf
wYSFlbrY+8RlwsJYP8T0D9fTkbiO5Day99p5iW6jKasWUe1QgEPsEcF8YGd0bsXJEuJxF7ca8cxV
5MzWtpyfji/TbdrgcYhjGILoFfpGY/e5RJrhWisrqWHjJsAGM/s0igECV/AM79n492f0DC4r78d9
6YbLcL6kWnAaRqJmOBcFhyf075VRkXADNHH5rMpZvrE6CE8PynfZxXZbJSsWe3glxI46e3dUDal1
phHk8+xctr7L1/rQY65XczgJlgW7JqGe/YawFiEZbMIAdYTkxL+8O2KjfL2Oe/Kd7/HVGte4holO
TYc/zNe+v9igy5Cmyc21zBP/H+7e8em0renmdjwaPu/mo7hw+hboW+YSUvhMV76pcNIOaLzgpg1o
Bxn8fxYd76BiWhvv7NuYa3J7K18fUinKBS84tE/lSMnKvXQHFdnxlpRyldlUOEIFMYZyWOZ83Nt9
79o72Pe9hshhhNI/XROURAvQjKj02fJP6df2yDbTO2nguZuNUZwRlxY7XB+KsX1F4fxe6Cwe0TWy
OcbyV8+cGAiW9L5QD4E3p4iNcOONdnQxWbBemeAcBDam+Ze4mmkXz1XlaND0ZT8rzRH30Uc9hw6j
TeJ1nS7LDY9a1buJVuiy41E595RgMd/34yuCUZ//qmzrtnanhYTck89Xc5MLiC0hBl9ISldRIznf
FXW19WUFwu6gixg9W/8YRvfsR2DlD1dRoAe/X01eCpJPr2kMU4LiXLmJoacZfsP2CvlP6Ahzr/XD
ziAGab6rEp7v8kPm2WAzDBy/u1PHs6FaaTpXUDEuR+tysYTc+JRLdY7gTbvwiFvXRglmcTHaLaq8
KKn9DTDFKC+j3Bo+j1/BeG2R7xEZoAFmI4S1s5vErYmdVODx1Yn+amYmpwlvnKpzE9/wjgFyYUZ+
w+AYulea7IJvSkJQEOVZcGnwv31m9eHxr4ibjSSYKjzhJV3atJ1Ew45SE/3RYiQqgb4Zp3sHfx4f
llcpofrdsDFbbUHstgCJgjRrC0DpyMYVU1a+S5zR1+S3L1nOVJOSIBQWMLqoGobA9paFeY/wemPV
AKVIQ9r4z/6BmWdbyFrD/xCUEjqENy209O/3x1q92pBqpPI0SVPS3hvQ6YCNhMeODtVnZ88gmdSI
7bQ/jKfM+PqZwhOgUkcUZgCYKtLOGkbqdsQ8E2ERlYGa1ouauWG+qJ+SXRwm/QkLXjBerzo0HMqo
ipmc3xeqPbL70pA7Vreu9xaZI3zNCZh2Yk26jInkis6tEm7gWKHAOtokHFOKLDuYHR+Yk5Hbfhsq
oSeT9U2R67gEVMaDA0KlC+WScES5iYEVkFrvlJz0d77GLJwNg9rdsp2HSyMLuWE3Eym+WrhUKYpH
hBwuLXIRYJl51gkP8qnb3nTQ2M7c1bQzDF0UuKl+mkCyYIzbyg3l9bof7ZzfA1L4JEX4goNeQ4ya
jAGZZJy+PXKVT/lB0yuPI0MhRVqh9W+cTr9e1ut+fpAtMiXnhKRBOEFgK4z+WlPdsxrMjLgIAmt7
mY6MvkqFcMzzbBQcuMPmj+UnQLuN1Dx42JWU3BL/XH/FjDCW8S/uzb3WcEY8qXOwIn+r1c/QdzIx
DGO17vretXuUpvUf+Nk27bNGVoQZ6GjpSp5GnzWRMbjQge+1xaDAGAeadQPVzebVY0Pg8hhGVQWD
ToSpSQR8yBO2fJ5WMO/W/qOy1Gbzu4AfmTp20VOVhmeGzEw9JoKyz3hXxDCtaAzwScYYQtU2ddQF
2sFInbJi+UkKZ83kXYekRNgYxDrqDx4tLoD6sIr93Tso1YYbRuqxlManq2y0ocRnriHIgtfzM1eK
kBQpOiu8IkFCCe5UWrH9yfSMffHsgxhLgCARbiUtbFU3BpJxjmbpL+/l4VWdzKqyj7ELZDz9zQwB
UwUC0w3rqH6YAdpHuFnngW7DNECPvMJ5Iy5nhmndRtV1jBbPrUvl7w1USwalYCloRlkHrsxqzBxo
bgJ0diWf+YvlGCD3TatxpVuGJLNnSvlv66N6ZlMufUTvqCz5TY5FtXagAtbQkQoSvmKMcfmvAFee
XLG/ug7ahzHd8R+uxnjkpw43fub4tryFaRZsYQGnK9lNz6HabZsixwY2zqB8NMdLftVs99Y2lif9
oZGclu+qRI5T2MrhpPJVf8I0g7JcKI1/FMtf0Ch6ffe7EDWiGg6GLjifobj0NbRa3Rr4/4YHJjh3
R1Bdb3ueBjlEdpgaSzajtnFtvPbYRJSRvHAyesdk7ECMFTxSB4BfpbQ9oNWJKMUXKuI+oj7eHdms
znXNKYYAmvnHsGzfhPCnqX0dn0EX3H36mUWkn0gI0upAa/bTDyTbEmQz3wJBLzMVEINV7b3RXL6o
tFvIRVSjlTo0YhA5eRUf/Fat1TmF1qhZVdt6Rwv1jzl1iUnKyNpA1kur59ep42xGdL/2CuKzbQqp
g3KFrzh9+rJ4qxr3Eq682ajoEzw72/YTP4xEYa0ZGnYQ8JCIUT6X/fvyo92xhvESZcCdY6oZCiCp
RuDIWJpe/2V/vwhvwv3IrUKSXK66OoNLqPfOvVanshuFGlt06kksrmA8Xw6mOHsT7RKkEAnhY0Hr
dQbXCpDXzERL+aBj9sCj2FpniaxhD5h7kt/68n9W05aluy52kcRoCqBi3yOSkTfLLL6zAXubpVop
acZwuAuScYw9bsLPYm4S/hOC4wcs3Ddx7Mo0IwPR3akhxSHup5fnsVwyriQAidNaLkHHKFVmq36C
a2dAz7JIdnpXkxsqDUjZjsynlGtn38BBGZcOQucrASOzqfAfeKNl3wVs8pt2y5VDHxPcCwqooowM
NZTl0EDPvembtCMLPU966jioSqLTk/jnsonZN72XHl+KdZOMw3deTYEsYbFSOQByGNMiznRSdtbr
lLiEhU834qUoSoSD7B8/MvASQMubbdxb1j5pIagDxB6qXkg/4VqsOvC6MMIjstEQ1DceOG+45cSS
/BImvWBngYO9rsJpBZpfAyAdXVWO/+nvGF6gngk1jcMxid48CORxStS7/SHCZ4tI4b4hl9JfOXbM
tXDM/H7bG46WmDHGj5XUg2mcC4AWyzQeRbD7Yhohl7jJNluECUNchv+1A2GrjGQvRe7LMxDXQx6d
FevBINuWQL0Ea/j8+dNNkwd+voK+pFpS3Q2uBKZWErpQ1HGDw3qlI3ONcRv63lOYQ09CiTfgyrks
bkMSg3pVDSpEQGFPs/9Q7/B0Qs9VNOwAMZXnGThb/8oal3EWkEgdytOjAGW9R81etwJFgcltOMpx
7MgSOxnmwV7pyW0mx2XHLlCgAC2C0dNAJz4/1NcgYPTiYFi6S2S3mp7SqRclK/FM+QKuOswDbloJ
rveKtyscJ6PDE2lK6ywRXeXw4LCc+8hJdTRNowAxGAFuVopfV2x/JR3hClFAxie+KmYoIYy6lWqh
UboyptZsDNVMz2RKJtMDHYf0GU4k6N93wHoPloLRUcAooyL1VXseSrkOoIuub27dnxKPfSVmnfVC
Awdt47WntHKotE9O5lMfkINXnkmgjdZhHeLm4Z5nQT7n7rtPWrkz191f+4kHaZqAwbBKaAUZverI
Gmil9kIJY8RZNGlGUJHfXXVbs4hWindJdZNTNHxYb/fGgN70LQJgH58GEtjxlSO6y49uF0NsucAa
W2W7EKj9kGJ2xC5ijbnQLCLHZG6PpsV9K2v4dxaLfkgnRoyNr8KmM4JiNpOFtI6OLMOFIk3ph6Mn
h7kvD6/ImNYk2BLZ1Y+cW9ctiQg88qOfUjli0ZIeemYrS8m1/ZOmoPnZCgdBrmIlL1SB6kTLVsrz
eMHUFhOJkoCEcATTvEivi+udwNRGUcfWVHKAZByjnsqg0ic25D1NV5086yKENvCEbDbt9moeieHd
JbRzUmo3V+0pDh1wdRCkuauA0a62+BxKr3GBXS9hMiSUWfMSnB3i0bT0uNwN86kVGpkyydgmySKs
f8ApnA5HJUgKvVnCV4TTiHUldsBNghW/6VqUmpoWpv+k65CgZ8nNx8NjPM8iqURH/aI/YBhFL/s9
0tbNUElwUiGPvb4BeEEdGnpEs/hVFIHhmIUhhiW4NAvR6wWTV1t5i5HpVUGTJbN7JYXg+C4rd8e8
6i3Clex7sEsQ9J92zwIbhrK6P9f7Y7X+Aovu4B+8XrLRtB/IGbgngb6FG/7bltVPjgEdvcYaYNNW
XXDFb9dCjH1l7GYGjd71hCjO6a8/TfNupX6P/d+ExBDCqV4mpMQoxZzd/G5bN73KG4+o4DIQe/K2
O5kc7zww9x3pijOxwuB3AJDgH/yFVKTE7IOsGAkCfMmvygHcfDLmG8bAhlzPLSY4csPUSntdoqKb
ermSxClk4C9hYHcvhiCOJyrvcimJqYd7sIN69/RDOMn/SBGenYkJxLmv4KfCfB8C3jisR/4n3jOy
SFKnpY1JC3HD09DbXX1idMj5t7EOl+plAfX6aZxLOqrJJi6od9QmAWxwdlLUvFr+TrotCZHOwH3Y
j0Vgc2FN59PAva1vpWajvRP+ySbTBpzqs6AIKnlXBUeeg2sT9G+Gfq+X9m+/v04re5VCuQXBlm/a
rDWvstmqamD+i35g9Pify/15sWkTvtnpktz1OwKR2RODFGVSRQRK5sXdzZo7COia3fCkVzGXSq4b
YOlPynI8rhnCaI7u0GfCvVYaIBwL0RCw7FS/MWDqQc+xmLPdreWtWLXF20XPmTbZf0l1mHVnIKSU
bw72n79GTkPPwPN8g4puQNCAx+wqIYgRtDx7rktfgtPCEN+kb/wK8zDhOAO6k5X24MCFhOf+FHUw
rFLcSHa8/TWMzab8bWCzondrq5Ucy5hl8F2QBCBu43u31kyHTPlMQbHf7QYbJa+mWIbu7rx7Pp39
TBaZjK43WmzuJpV+UR7cBlrvwbyqm8ZEetNTcOejfQD0cb+rEbYP5k+aV6RaeS98qsT6D+TG1LZg
ROIlfXP4g3eYoTGAnq+5LEeBn8p/FVIKb3H6tdQPcWpWQx3BYeMcv3wSkjc8lAiaqENqdIsMwEJk
6pr2WxMHyBQQSz09sa1xz/ombYvnkVVSugsrHWPvdXs640x0fUWp07HJPHlDZkmS+yifgcV6qVCq
k7pFkfWcfwmLzQzmskvdmG1kuEKdXzEe9NLCTaHTeFg7fVz32GERh6/MUdU7YixgyJ6MWb1tgC0S
CIRUmXwN/i9Yf8yyZbgKzRt7GUiFp0WZO7ytNU8pdoYRPRl9hc/tzdanO3FHnmuSP3mwaS0CBLDV
4ipCcsbDXYS48ggnaCm6odHQNj02frJWunQAt3tdtLCnBsf5KvdEZj/3gbn0XGchyRo8fZRQ+QfL
mQWOs6XfUnAiSKUWunRz7su5hqQqiTWxw2asHeBosA4kDxJMOeoFFlS4QnmIycuYF7nou81es2NX
NqAVOxcsmb7dDEH1eH0XQqj16cGN2J8FOI/Et2qss4kb9zXzp3c8uSH0ZOiMdGEawMjWVBSPVuql
RAQRWUThHsSyRNDDZkWSaoKgoDNwzpFYr7tPpsyH0tnwT9s5Mwor+Kjke6s9vkKji0/1n0fOsrbr
3+efA1POE98vOSkJlzID1ONkb/G+FSyMC2zqkjHiIQf0YqpTyqUHsy9stn4wNjjS35eTFI441OnX
f1dFEFvJRCNZ92GvNjGDHjmEiQ6jPwTSvA6I6p3dOaWWKIwj/zGTtayD+lBKOLhj4j4RUffhIi4T
15ZXVsO2zu/z5ynG6Lf57MDpIfKXxFigSpqBWmBfxNbY0MJYh30r2rxPXpWLMRB9onldWyAdwRQs
/mHIENBiqFF1r1Y4NNeksPWuIalBH6Pj4xiKgZN7fhIebZFJsoooXmzjl0iZ18F1sbF5LsuLOcM9
7J408B34eb5KCYybfLzVZ5jxc4MCLXiMcLjsyBDirmej9mVtY6kh561OhsU2r/Stftr7kW3UXJwD
Gxks6HmhM/+VkiwtE5bGckVlzX/arzi0ZxWgNqm7pF1GZHiGkR79xxak3N0COPuymd6TaQwY1W1A
M1B5MqUtumKE43RcN0DSziwdSjCpB4PmhrBxpDIwUncmewFg6mrzd01wo2k9JVlT1V7G0tE4lipj
4bzjcBPHiDdC8UJgbBMYf61995qAfLOp1Uy2Xsv5hz2kQnN8A0VniTj8t6L6iI0dWuUVGzTXuaLk
reQokxWa0Blso5C5girKvkCsqdY7Uy7dQsW8pQybXCGHE/fTzdFOXofs7Pj3ZGsUC9+2MLCVaBBy
ywoyIy5ycFce+J5XJd6bPvySLJjAO9OiupjtWMuLEaQkuMJefdWPeRFkDET6JbLdOSP1Ykt0YPat
kfoQlwUdUC6/bFMANHO+dT2VDOVMu3LQpGlXr1+dUcldse8llQ4XBoFm7gvHuRqVhjN+XMci0+2N
hJR7yiEErlhR0EvdCbkJfDjpPFHwJkoOvqer2dGUntbjMM2Nck5oXoShP+dsRJTOxTY+nDC422nM
KRngiFVwXc9aiHCzqt183uCouQ+5GRSnZQvusiJsnILz/fnKMm3Eky/ROq7W3p+jKrtnQJ5ndyLp
eVBoCha9mpM1rlCEaLR11OYBSRxIDmaKs2JkT2D3fAVobvYzo+39eG20BHZbycU3LSNLC0C2HuLY
e6DUMIt5Rgm37W35qJgJjby4sq3qJ0dAShhrpeECRnymP1uPcMNNccXrqjpXIgW7roArukCOSqGS
K0Nh5XXTIbA8JXZ8x4OK/ZvkmuFWusW1SWa+Dnx1Kd32OcwVa6MlPbomkIQs4GFhdF1BT0Z/RGcD
9LVKyuXFoykP44LIN46mSJaO2XZckA2lnhD5/RovdKUdqr+Hzz5LBU+C2lTMNU12J3ic4Yf/rTos
KA0+xAgkpnvZ5D5plgzzBSPxTLHR6Tc3Bqx0c5FlxFRCapH0l5/rKGMsOvEsyfSZzqVNDsNrNuoG
oQQ6+9eYWqDls4yC7kAWHhOAahiM/1y8Zw20DxWj2NfR4Vpb/R3Vs6BIuybrK5JHHMalLj4FFbRe
1u2bXjGlGE8wh5N9saScFREZD9mr5pKQ5lbkMWUahM1DoRW7+VZVYhWmx4sxJXMHeJQboydDeUak
U62M6NnlK894PPKKrQGGjdk3t00bn7SIhZB0V5trR1E5ANMCHc9IexWRuIeDk2zV4w5uGXYk5w7m
Se23dyfElN6OB+r24tyyebRLT2AytxuLH6FYQVYWiNFQ08pQdyS9VS+ReuhgVU4eoUYy7Qek2Quk
ROxPgCfte4JLb1QLcVJJw4s6vF0FeY4ZvmmeHX/j8sQgFdZDFu11IyS7rB2tdFxQO8Swp0CLkAuK
YVflNB7DBHWd4/FHXhdxBbeZkJVYy3fp61uUgiTuTxhkcWOMmERwtIRwHg93aV/tXKS7LxsePvVz
G3KBUVZEbZo7cjZHDenmGTEY/F4yhrvhOW4I7thcI38nL7+uYAfOabNloC7csGP88c20XFPKKdCY
1OfUaeP/Oo4zEKL4ZIUCz1uiSxvvnFNWm57AGosrXMPoQUg2RcKgsm83mQrZ0hqyauHA9ijElaMu
lCrU8xoKWiekUUIBDQjTv40N32MmrjuUVFqcghHiqoZr6nchHw0+SBogDiKw4nSMkTHRNRZOS8zX
aObrNZ+Oc0GnET95Bv/DJ0ju4s7PMccISVV6ro9WhyXUXVB00QpN8tZW4NddRrqweO6re8r2wFcR
qY3UpEgfBQfFxTm3DWFnzDk/RUweJdSZ/rQ/IuQfYOgjksbEvEoNN4SIXqTswbiAoQlTEr8en8wT
yMdvP7MzMW1eRDpNJetIstW7Zqcrr0bhQoyhOtt30iu6Rhg1vFQWK2RZhecX/Wb04VsXAAVM7vKS
zHvpdKGKSi5vP/tSa5I0qFIdwaSl5KoarC3m9HJho/UW3umD7Qu8euM3N/l7ffLWSb/CcOiGyuXX
7bUIrPH4plvNYnn0XD6MlaV+2Yp9i2ChBfSkVo5D60LF9VD7ZKvYGftkSxePGggn9fnyQIja8L22
uHlcVykjBLyhQt8nVoAF1lmb9+16ttPuO8uEvvdCe+Lztzgh2gzHvSJRxkIGyz5gtndyFtDh4XlR
G70klkuQ9Z7I9R3xnnuKY75WvRFlcnf0GZdj005cAYzp+okYD0w+XbkjITkJkVNFJYjch4zMyrgV
3AIx40tRdaDwWAH5BnX4avBGEkZ5+ybMmDCdvUxlXpvvN+lR3r+41DqvWwj2YnVuY+GDPOYzypbU
9N4t+bbB9SxlGDLAXssnqflsVooVg7QnZf2CKURPrbf0H7QpGt5PArXrX2PFyjDg+edY09H8U1M+
aP8JwW1n4jSt8A5/KpoTl9Mzcp+Mv0i91Nt6JWAMsWv0dkXbWkrvxO9q6+nlCZttEFtz+IoHpi7a
DMZtEEs5rE34AGSKHiI1ZUem5Ugjkg19iTu/RqLyBCBp1DHyN52N/lhnMPIv3zLEucOywcjWwpDB
khGbtJ+rnRNJJVt+TrsLn1cSZDysQO4VniQRhCMngnzDPQCIE8KDGEJog2+yQomb684uOG1oo1h0
ep2aC7gYbadVY+0Xy5Fobyi9LgSvpd0w/LKRzL8smHxLCGajSEzJrFdUvdWilee0HjpSWpNpGn5Y
Q/8nKwe30reAu+6DLJ2Mwr4oiOXyfIqNiFK5gxIAIqaUZPJNdnfsUgdCFSGWbOwKuRlqI6YOgEom
04AnBkoH8TIj95yFetXsJvr8ZCc+KAGxq9R2L5rdc8HsRYrRISMENMKJyKFIg1vjVF2ljdXiV8wR
kqqjR0AbGsu5FW0fhYVndZqdMgV8kTR3IbxNsaZl4anUi0Laz079E1Awc06Z/ao0ApOACd7or7hU
tqQbml9PeBK+lXKxCrW5dOuPmLm5CArGvjk6FTMtDMH4TD1yyFAOtBVBWDhH5Xhlh//HG3jO85kc
KWYgUWko1IOXYKZ+TPpDPaz7lMA1Xo9aDXP11uuu0sxcRlbH53tzJ5UjLs2Y4WUhQp1S9urP15uu
D8ThkFnWxjX+RzaBY7vTZjtl9/AGaN2P2BjskitU502eiEWPiMF9VCfKCnBMQk58bn9ik+IvEkSt
UClJxTNQH8/BA4whlnzdwmg9yec5rI7Glxyqn6krEiAV0/XAJxjM1Sm6tFgUuW6HHZs1ymZ8iq07
VtHEbsz+3JZh3ECcIEb/mEKZjL83RVlbFpZ+01XaEmmcu/Bc5jNNSwdF3ix2/sP2fB4IIXpIfZHf
F0znPwT/s+4l9TI0J+K2lzUDR+QFE6NpJkcpl5QyOJ4YEbqOvpDsJMhwsxtPKPuwh6PKJkzJInSn
hpX9iMNxGXwSiGVpFbbfEafPuMTYeOGC++SVFK8zO0/D1DzRTVwHOKDXfIXWIokt9yJIjrTIs8QZ
XPdMUi8GiCT+Bi8/OArV9kP9D5riXEBlA0Z6OOcfeH+FE3fObp5vmjs0WkY9tOpF1OQUTMTyIM6K
ETuTkCQltC53oAlzUPn2EXJsFQl8iN88lpeLlQn3aW8ZhoO0FKcjjJ4FqOpSr7HG/njoio/6DlgB
RdZbCm1Id9sOIdLaeC1kMQtdXxMMw6+DUe3hHmRpD7gO2ArsNuahO2b23oJmILbvZnJr+7DNq3Zf
O6/MI30G6yQggxLxMU4GGBCkeViUHZe5J8eGqGym3kirhMX2Ps1mMjqWUY7MFxuFVe7qoDMCDldD
m7bYNWEopeNTPyVxOP2jGUyyr5WuJHVIIfUxmZoZtpT3XEu4zwEAcIuEMoFy0kMEj+YeGq2KqO84
WVY5MrQKWFVmVyADUceDBYkDqkU+IkjeFucQMpYem91cprraLcqgOeo95j2UqUnBvzjtdvwnAOmV
05WmfmkSiAEOfIxbx6bPhti2oiNgfpQPmzgtZnEXA6idpgU88HEphYZ5qXiPl14DXWs2Xr2xvtaM
FT7TG8K79KcHOrQO1sba8pA1EdrkhWmF+5F+UfCnY6wie/g8ar223IeeJ6BOUc1Nx8TWeVPjn1tb
B31Cy+WYIfMZKrRDuby25AQHjcBzH+8Nwg/uq7BZu6JoHjs8CKWzzST+wyUXAGpnF/L2rlewplpu
JuDLvcKOemA0cv26n8p4aWshBZtzhBEIBL8GFLaIMDJ19jO32M33VpUZBAN8tdGeslO3AsaaekKI
oKuFwiQHkbtJRyj/vyccZ0dfDAgLmPyFiSvXnc9hqIRbuHnvvrP/5bG6Xq9OFoKUGm+lAo2Ipk6z
RjwBcfSiftH1tCV3A3BBAdWSawDftOM0/BPMcLb/dk7LgZL7l/DMSi0rGpE6inEK/4O9FTPYfi9S
pCmjvixCswAYxMOPsS3Vki1zkHfC2KBa66bavN54zynftWV3/tsyOxrP6OsYCAA2wJMsZZJW7uRE
YlGUS8vQoBWnr0bHDqm2n2cWod39IoA8cFOc1ZPu/w9BokX15Rrxb/jL7sjB0d0iGKC/sJRLKUVE
XU8wnulD1qqZ2g/a2C4g1JlJfOWw1aW9PhaW7ZIVj0y6x7G9mO2btVJj1/fAgzOOh79NxUztT9rW
v/d2Z3yEHclErj7sB25vzmhW62F6lqoZPrlL0GnDipvptcDMMm3q1S8mnQzovG8N/T++EDEdV5ly
+lyW7wd6qea2pu+2jAZrH8OnPKkxqnnbe1xTHFncdCBfltn9lNsJEFn7egOzVmuV9HTHlDgVw18k
MXsN7B8MQWw4w5Fep+v8z45zXD6JbFg65j0c062nbmJFyG5DSKe9jqkM0t7Eza30SARC6o4/bX9R
Yls9ZJ3oqrhFxB3um4w9ucr1MHcg8/9K5UuCFhSBkWidg/s3fEA+vtMpU5RtjBk7NdSnxr8G/9be
PObM1TFo5301so6Qx47FvilQelEVdUwr5XAsmzlNhfjAzeIUU/k/OXViqzK5tGkZzbNK4GVpRVQu
bf69yiZKgRB/6/m7+U/AoXODwOvkrDtML+sPddwVsnyAYJvJFXBskj7rfylOSZMfDFsOtN6qf2ln
cVjzacfT1G53+FENysnEroNxSmeztZhJWzOMM7CkB4rXTNhtVvT1w4EWn1kSINJd/j/NSwEdTtXd
7AzvPIB8GHvQNN7xD4aXG1GnQGmZ59/XNwk8yabr9bZEQL+bu4Xihsk+fxCIEkGeQqTnEyISkZ1O
wJKx4V+Ehkc2lX2MwEhAwB03b3YEvwVDTj/MlVzwBqH9aqI1nmL3TQIJ4EqcjAPA1yanbE8Pnr8n
/jjVv9EXwoMuJsvLK5GfzeaTS4T22ze9xhySrUbwAP2uH+71AzZkW/XsxqxzaQn1wQRb/3mbfC8x
3HArXhIGqbItbdVi/QE/MSn25XExPL+Dh8R60YaMQzeZM0KwSyYfmxFaeCrrtUjgf4L18XS3w7ey
8oh4kvODV28iaC/iALEJNc8vnYgSclkGPmgAt/aiI2WGs4+DzORGtYVq8pIkakT7tUJRpzvsIqgl
G46AHFAWdsHQiRpUWeQ1XLYs9koU1D2y/edt+5R5ZJFVd89KUfAEEo4omHSMCjMuLGRWpTNDsnUC
iGhB1F/xftTiIFMiPc7HIlw2/zeHoeDhyZ1z6eML7oqdsEjnhGI2NjMdzrdcGiCW+0ie1GYYxPEW
P+VqUHZeKH2TCc9pZcqB2N8sUemwDR0QIlHZaCwhybtSnxGMkYFZCGQGd1kAIN8FWpkR5GgeOzLO
kWEHG8Tp5YQLbtxWJqhK9XjCpLAhwq/GXvG7nFoLJaSdKO8UyBnNKR0MTxtWCN/IovrUulG7zwFV
7ejtUDw39gx5NHjL/yD2hmq1PgufWYGajOVIF7pVau3lcu+OLq1MRGmgTRxJSSdyHl589mFyRBrv
0qHXZQ6A9H8i1yFtWBSEFtvJj44ukGN1ZZqXkDdU4lClaRP7e0YlrauKBwwg43ONCQJIkEOqAbC6
z4jKbLPhoRUC4gEpDq73LRON1xfGQEvav6WzgbEf0zPIv5bNzwqIzfarYNnvxc7FGMQCJqGwq3oG
vDyzFredeZEUXZtwsOE4imk0/+1bofjVR8eqBYqbbRROvSxdL+LJl3f7XMb3eabswYZINjVpzKbB
45jNKz4s9gELMckCyLIhEZJvQQs45EwRF72NcKld1grhnSeC3a1fRFJ8YoD5hBhck48irBHzWNUU
yX7/Vv0aT7VrMSexLr4FcepPA9walF/G9JWZloFpcg9VVIpwYU2AaBvNfCdEupmptrcTPjwGk4Lt
dF7hp/FcKU3JNSOjfkHCYTFE4+/obNMyRyre1maxehrbGRjoLXjO9TWTkkzDzu6Z7/i5tlrkVOGa
MGcvU2sK+ccg0VTrbGOtM03AEAGDY7fE9DPi3/U6Pq1Y3y0xpkUGjfNG4rkXQEFqsqRdWgvC4R+/
SuBs48pVQIDaWDie1Yvw94nzkwqsmM4OtZ/FbnqaORge9ijW+14tccZlj2rsgYKlu5nuB8GAesuk
qabkdjckdWTOKy+t2tsTiC2QQiTIy7jogr2s1iLqr8BHpAaM1nDmkWJuzc0p4lw+GADi6dwNUS42
XAoX6Lcmrpo2g9KYe6Jjnenpabq3IBCE8TF1sd+oT+Nj5bDfGUvJPvrgMOyz5JJEsJyVG9z3AW69
NelDu+47wuE8ZlrcbkcMEaLc7zGo0KNw8OlppKH7kHypjTCkQ3vIAorSfnlDOz0jDPRtWO3h6Ksh
e/EOLSWT8Ixd3KpU2oDn6+O6ANQqQUqxcXBYX9pVv+zzx3K/q0eM0tA7chhkHM1VFh0Wkei+cv8p
m5ZRWprkS40O0bxMQRXiKW7vJyNyOTUhXoDO6OSUwNOYBRVKOaz8z4hdDdDKz0Fu6h+XKrlg51mt
SmzC5tGO7RelrDLNNFbBWMXl98iI+GT+FqBC/6SkfqS3mm3t1KjTb3o7PE+3zKp/mgREv9ZeWnMq
0Mm13Tdbg1sfUAjHiYcyEh7covhP6DJzjJm2mWRKMHDiMYdV/cvJQ1bUpO6aSc1HjB9ra5IQWvDA
wXUFHGQgAbmipz7HnkhcFGGHtIMXaaWAASjskQ0Vf4dXMx+qW9i2471f6TD7XvDKJPevRFkAJ0Nb
B2CkKSEtctMG/HgjdHxUKaMd4wsjgCUxueihsrQ+ASuZxUg7Sl3CtywJb6Kr6S/TNEBGzG2bq6cR
/eOQb4Bv2W7BzrfNnCDAK1Try666XcUEVFGRoDPLN5y0xgz/fmMiJzPOLSrvLk8lbzwsgpGxQ9KG
P/TzXopOvz0NgVsvbDU23gw0AqRcITyXpA309/lj0F0K2MeAkziHoCmNsHIwEOtBa2kOwPoxzPQt
jMQzoT7w6rMsX0DhjOW4g9yNGbtnkApmDA+KUXZqp8RPnyFLA1EXLmZfRLw8ScqTVcL9VXPng5cb
ajAqT5Io1Y3CDeVyhOPzztACT2VX0ytgy5S8F1t6jr0SN8N8A9Sedavta23kEI1kixPbZQpg4Vlf
Kca2L4/gPRu2Vp0EObWe5Mp2rNqIVCt0BQKU1icrIXmg2/ei7QEDA4V2Rhsut972jA/lqJjgbXSu
WEPQ8DmGsbFkwXGRT9TS0WGdzvAdP8YntRFj/pmZZpDRMia2wA2aR+1yHV2cYp9o9LdVMzUQeH2V
jogxgoShaguV/Qa0fOn8gAvoubleZlj0dR1DXEEkirHmAFUiwEsZI6gy5MJOSSrU3xZBS7do3CZD
tcWbI4yscBPPo3ZPvO/0BfTUhjckcfXAByn4mtjvrlWEte5gMkHeJSueDmokxPNWo05HYlPwmNCQ
frec7gm63aMEoQ60coqwz/OO1KbTRG4CKrKTxWkQ2k+J18AV0vj50IRawADI8JW1jde9DGpWcqFa
CSdu1K77k5z572dnBzbtYLIsptyuA030TKVmYEDGE21gvRXyA4bjDqcUY8slKKLXVV+TlQtfca2i
npNjf2GDWfebz6LQ6NeVgPvgENqUErCtDQnif8qFBGO9Nhq93rPRhVmkFVMGMmtT2z9n4WMbVU86
HrFclWVlHmUBFBQ8bebgQzEXDFx14mvX6TxwbbVSwHQ2L77IZCfw3tHixxgzYgxFvkeOyhn81pRJ
mKlo6SIHAw27s6Pses52Rjho9FLd1sBaFATL+YHzTVIyYWxq60BdIyk3VpEnnNjpqfuSWnPONJaS
EzFSIbt7xU1H9fTB/MXHl1vZLYs3kUYQEOG8xzzF+S5Vv9CqkD2hd7U+/00cj6GjT4qiDTbQpd2s
6YMyTwYvFEvsuzyUjNWM63e3RpQDd5H9lFUQ3u5l/TPB5pRO0N+aylINqxNwTSKO4Bs+V04TnES+
cKjjXwhVf+jstcHlks+b+vk5aHoO2iiKI57CMgxWJt3VLNH2n8vszLX2/0acvoXBPHSYPU2MCHV0
xX4KygkjdCSxHzPCKB4skw+PjLa+g+XKdde37w4kbk1YVwWAK0bVjPUPYiIpzD4s8VkxWE04WF0A
TiWwRuLp0uBWG6JUtDEljXU5ctQxo4LWveBG/gj/qNgP6Ln7TD+2s9cbQ4PJZRkwBwYTpxH7LtW6
BIP2svA5TcJAEydbMqaJsrTCdXlIjee/AHQ3M8DtAguUG3/Km6znKoNvToJ1DumCSZIc8pWTO5v2
1QRjVxrgq4OY4m/gU+psK4rH/RC3wdBl3EreZwcRibifMDS4MBJEhC7zm50Q8n3EXcsYg7F8cEXG
kMTy4l0V7xxja2/cPdReuANQVASWykxHyE4mXuUtIMiC2kv/g1hfWpbMlkSVlNBh8oou7Dsq2OC7
3v6rl4vQCH6cAFYibOgD6///G2mHi9T77n0AsKHIwd39tyVBmPknF62acONP2O8LnyByHWGHrN/1
p19Yrha/uqrz2b7FZgp+7zPJrgDFnY3K7jensrFlqgLRYYRRViHyCawd1FZt5PTdTHodZVnmpvDA
BxdjZQaImnC+N2IrvFFQUEmO2AEZgOQQ7kqp5O41hXz7q+xfKf5jg/Ui/fjdsKlt56XAinKwUet2
4Ejw62H+LMV3uUYX8b0KCUSXpxLfNzLJ56YB/MjeWDmtm9NOkKt2fhsd9KqfoIQYp2GK8jd0cgHm
hLkAniZRZzVgLN+7jCb8zxeh5+cfHr3IfnCUQqzDXpopAhk1z+jbHQU2nJGXCQuhY4ULxanK/XFh
cx/1D3ZOYRJ/A9yWm0ThGMPb0JkweAo/+I1zqvR3O7A0M0XnmlQA4VYacLpo85LMRMFCPefSDbDK
3TV3Pmx4UBYkou50VRiGCWdK383zxXQuHJPMaGJrYofrwKjqWd4asqVpgrT8ZIBbMlU6KewtCBaJ
zNxD8ynoKHSBtn6bQkwfx4fFOBU9F8pQRYL5pXSPucPJA0YJjRsxnm1ZR88q93yXznE8oo9WGtoB
fTg1CvGlehgeuDb68t2YZkmnB62n23efnJgzXO1vBrHAqTKjswDthWG4ybawlU1o+u8pmpSvSJ0X
PI78BQ44Ct4tJcTuT5nNgelXZupCdsmD6a9J9pFHJci+QWR376UIOYmvtgONmQUHRH8c5VMO4+r/
qxD2PpUvD7LGZz7xSBVrq1nhH6l7otNUIXNjTRPI6G9YOGZlyr9pojt2TGefwrVfaNAPIYb0kr1b
guh76vDOuXW/F6tXOd1SO0FL287xWn3Qp6fmT3d1A2r8AM3+JNySL0PmH54HQvvG6ispGdLswssr
lbu+4WghnF/0abZXwpDKQcKq832TJ8Kms4V+oJuWyuw8mQPpeQZDheH4xzhJZMEqEitAT5ZlbkKU
a/35UWTDPQkpMp8GRDBniVkLUzZ7NwCtMCyUFJM/JBpG9Hn/lYHVm4pZW7kEdGrtY4uFBJ8mfnSj
jpwhSJqEIb5ZBydbTetlHi8iKr9HWyEGsOwUU/dRInsrn0/88hw2M/JQU5Q9lJV44z0EodfpEZju
d6Zj1FcmtLwX263iwIXAhaLPAUyRtahoBW6E2h5g7A2ay9WxxwSshRH7G/uH5GiuM8B0bRZBjBCC
hEztkG8OW8Q1hEA5Wy7l+FhfQkyOW6IYNlYqz5YAYWkgvKIacfrSsTT/uU5IR15ukfe2Qf1Qfplh
A6NBuH7MYw5Je1gmAsbFWTTQAD/9mCe8Sunf5r9px3If92f9Xvd64xFeQcTymmg1H4e6u7YqBF9X
2OOHa1CWUtlQy+zUbi+2EwZrKJRJ0AQkCpUaHSMSQfGzMHndD/N0PmT17x5xv20l1u4fDFXIrAJh
DEOsJsvMdnXbzs5e9pB1e2lfSvjcNPsaDQUBuofig3lEyXAsXTMKrAsHl14N8kyv81nHKSW0nJem
fkS7ZAeoTNdeVYyGEMfUgv6suACUWCr8QRqFIUIyDeH0XJOhbXHEU4PcEpe2vZz31cGvFI7D2XAO
DuTeZjY5nsgo/PFOcsQcD8X4MIllojvuZQii0jh3ScUUEFqOagkA/TNFC7KnkCN+9Bh/0AViN4fm
gDW9jK0PU1ZFi9bcCo0e7oZN5Xbwi7ogTkBkZXg6XSpJ3DD38X0B3yVEbLV+iyHLCCYlesRs3YmI
VLqFwA5OC/chw1MX3puS4VMOAB8u4PZUvtgjF/H4/3qBTu9WzfEiMcu7muH4vJLdkEGxOOJqvLOr
igpMoE1f3/FVm2AQ2ZxX4kIAb99/zJc9U+kSzM7KiOw+hybUFGn6CIaWMckxPg6jnrjRfT/AULtj
LjwrZx1HSYkuEP4gLGfhxrkMRLQ8mOITcOFZlkr/KRGPTx2vSpKjaugd+OlAGHUiqvwvWKL2zTwm
/9giS8cZBp/FPCYe5A5W0xbaSvxO5aAH5/mciDDJcJQXMFh3T69Flwp0dWIXAsZE6+c5R2jgxf0M
VoYrWW7d+x9vVgZgx9cGj7j55KpM5Fzb7HndqTPN2wfItVmQPEsvdurvrMv4oAZpBA+TuWDG5rQx
GVww/avCnGaIGlNv5r9w+CMHqTP8YzP9i1XFObB+wAA7a1wWSGAcUMMrKS+bSZbunylnI0YPMpGa
etFvW+ZqWf4jXd9hs3eEoWKnlYU7l/pXfzxIQ+/fuxb1H3Fo0MobRbi1Z7U3yjSmLhxyZnKaqunk
EcMjQLTFYFOooBPlMeTnSQbjR3sp2U3OFCL3c0gqcpSR9WZQWD5gmlM5RhRU/eQ525Zy7EPud7RB
Sf5SHQksaxSAxkOhGe9w5vWB2+kDt/LngcLzrUDMg92imLI4bs2T+0wI/HJhFqL2TxfCgrFWxzoT
pnSjftZzM9cBRz9RYsVTwyPAQYLl54lYB09ItEeGzMGq33EB/aI4vz4gTqHB4wawb7Gx/36CpaUb
YQiooZ89Zj2BRpQDmKLXgXCBDXR+HDuioSsadzs7REJ8YdgoDKEjwe677BMqz0n2jxjVoVaqq1du
RFnVEddYXkldGgEkTOldRRxWSkDJANbDcG/cu7iWFlh9MvMJMmkUoZtLKj2EvqYBb/SgQARCWuzE
B4DnrPJFtq7rSxFBv/lQOGB8ZnX5FLjV1UROPtJ/A/qgcpc5NJyR/hf7mHe+pdEgcT3ImG05ZISN
eGXu7CFRYTKIGzHAjXeIlPURLo0JX3q2kB54eXewsaAJXIxCJ4Hp4KzlflSH+yqlYxqmMX83Rwub
RlerI5o1wqjPCv340pMvYVN/iZn7Uj1h1b+7qfm6YxruJizMoYcT5cvberIZZvNHg2S4o5jrY8Jh
e0YT2n8s13um0BbZXSQMFy24p6axCCAFx/Hy89IRVhjhUwXYIYwYB3ziHtDtgIgzUt3x24mYQQSH
k0eb28vgdbEMfY/uh18hH2lu2Cdu0mmvGgbOPSPYMwAFozdbX1iNUGyIeFB+2+nwWFdkid3Q5xkN
Ln6MaqOSX9Ed8Dwys7gDzzLyQG5lEQiRl5z1Hef5QAX9M4245QbNJeQAtoOSDrXZP0NcIBrl8BEQ
pybTQ3OkP73TR4TzSpPg3TcaRb0mNHTXE6iFJx6sSuwECtqMXj3svXCxlK4eKWsSl3VYLou56VOl
DRJBLlrJrrNKoTdP+AdVmA7JSHymD2PVBgtLeBhGPuDUnEQ+wjpqhQcHxQuwXDbQDHKg8/X1xaDd
Vfq0HCoQD7rjHLXDOC+Gg53jdxhpFPZHIHpA26IzoCd1uMULOYdKbDkbCRuLNenRgJo2qR9Hz4Iq
1vl5EpF5QohJULh+FBU45QV2NEyj0chcN9s0aBMfCs4EsJ+d2XKrl81whR4vZtSxXmz/RWMWrqmF
WbCNkvwIBj6LPrTMbMxoHMreymdoS7vf/pah10RkSkdt8foNBzp46p8vBzqrgB132+HPPq73A0hq
8baGDG0OR3/BTL2CRsgeK3Vv7/oUIVHQD8BddAypHDVQF21jlA13hhJl4w1aiiwtA8J5HraKyBDa
tCHHyBXCE5X6OUuMfodehmJRATNFrr12Jufccz7R0SagMtkreADByw1byr7NKqpbyQu8aXq0NDmq
OZqOI0zBBwEwwEH+bM1A/lioon3gKF0lQ1OKoduN2P2aYsCQ+JXAg5VTOYCBtg+rl79vDf2crkHC
+VZ9ENlGiL5hW4pLwMHr0U1KuocQYxcOfvqYGwOgDNNgo79IoJ4Qr2CqvxxGs8yB/khR6BYoM/Cj
rAPNCt+9Vyy4KKbjWkn0ZIXNV7l0YMyBbhdt5YjW0aQu3z11Npx3vg4kybaveg3cnx1puf4dfr8o
M1Zdo+vvtjGkdubID04VUKNTZjNMMOhEksfxyczGQRGzLg17yX1SiSe4dcHknfrvkYbUO/nYGGGD
g5e6kJhWfT1C9SekgGhI+NWfx2RViAF0IQPzbb3MytKZEm8K62uZaE7ygwRd7T3a8U38Sxm84gUF
vp8/N5WZQegjLDEASjA7Z8QA5lnYMH2zlG7cCTTzNeI8uY25bvd3GWCqtUYa3ymIWE9sq8POQpfU
EwgDCo7dzbwROzgLQ8d9lXVwuHTwLttbmjkNorgbBRaa0wK0L4VRz+L2PD7ZYaVSergChdSzLZGj
WWof0M2yN/j7tm53o02FtAqQn3MtUjzjCKWQPoE+nG3FL5vfsEwcJOJ2Qx7D0LQYMTlT94nGiiRX
CN3bWiGRoWdDy6/XLplxHfsV8yIKyXssB5d/KrSmiIAK9f+Jb263QWDiYQouS8UCo3EYrpTlxbMn
YnOwXygMcPzwA1AXnEdD0CregvhY93kHnJg3yDH8mJq+yijKTAcXcEXkdklxBWIlqjozoPeNrSmv
8/cJj77EiLBLHHKjVeVMWjgVUpgg+11Dhx9rzhfWv66f0TqPZFHwqQAm7+GzzVd+boMn9zZiyGZO
DCuA8kyj0fJ17/808vDkPwvCrQEiqUGNkoy3v/LgNaQ6h6SaKA9XkDtZWjdLCpf3D8fPijgmQZlv
a4N4pgw+XN6ZSOc5Q4iQCmTxiZoyUlD/+mLvTsGqJkg7y5V5D5HpHlps2wtgcvcaRw7m7Zo7UJSD
yqAT4CIrOqg21BZLSjtp06jsBVlG2Q6qjtH12BhOnlaeH43h+QmbVEoqAEoRugbtVbGzQNvFVNBH
xSZXGE0u1Ncx198+DMOnpeU7ufdtzLGySxHi5GYlfLX82y0sqmbxT0hPYV6XSAvgg3IIbK6MN9wD
2TIW3EW7IbpU0bcJN7u7twXvIrxMuGkbZAa+LttH+Bh8xzEour+9xJ1C2IPno3ZFAs9DZoF5Nbbi
i3rcNa7lBXQJZRIyrH6AiMw4IZY//q056fUggfTLoIsFu0UgVPPA0G/MPES6kCiXP6Dl7hx/zhcn
8v3RNdIYqtZVvkeC6z0+rTvxDXpCUMgAmxnpZdIt5hBDS6qIFtGA9Q5489A9BN0L6apb/qeQZhWy
+ULxvv9oaJzSE3kbcJA6EyPpdvEeM0isWPsuMzaoo24v3V6uPTz8wU+4451FGDrJjoGxUKzNo2Wf
Bf7wpVKumKw77GJpTrTZK71C8OqyGL5a0qKJmSYKW3/k2i3KmrjcX7VY55RlDikDHEezkWaEuWv7
S3CZvYtgslwTPvHrfJiLH0EcRTWDG/Rp/dHgwSrBoc60dX0I2ZvQeanbtb/E6FCXLtH+ijtFCbNJ
wZwGb3uVTBpD+TdeUWYYSrK7nyjdSNnDsuxExWh/PlQhlBP9fL4nIrp3n1sPxOVoQGuL455LiOD6
yp6C+dHvvszMFETUDdmZp77sL6EPiIYOcajkvSfMrfl/gUKptTNnLtQUn7i/teEZXWs+SmhfgYZN
lNEGOwx2v679QkTu9K8SDXIfp8v6NPRmyTu0xwIecnqlO3ty20h7n7rn6uA2IoAk1i8Pd8RuoQKo
ff6EKdFkPtbqlYYmaYxKJwEsFhCQWWOJD3PR+wgQDNZyv5RdSkxJdshZA91B1WI1S+RymvWSpT8k
+jxI2UzezXfgCUAAO6Vth4PSF/6cAW78iwDGx2nrKh9p3RZc75fnbWcg9zct1X7tEO9UXKjfUgI6
OG8LHO4zdEBHM9UH6p3k1JOivvvH9sglFUnGDm6mNS5nLiD8ixN2vPNYl21s0SnpukMBf/y5FS48
IlH0OmjDdW7n4hrBi4KCWCG74H6qkmhXFVOozVcwciYp6Gt85VO8NBIM3ucgDvbwi71swLtucTFx
SOejYM6GzfJvzO5tadVvKm3EeKJu4m2ELSaV3kW2VDdT+G/XcG1s6gOBtqzWvnXgZB8WQQwkU+JJ
UBmsvN8zhDBIXcNDnPP71LdcFIFzPlLZAVVPmV+QKyuttoj6GgKcthvty57gZ5KvKYZtaw7MMSL7
ssVouVK42f6Yi1X5X3ssLeB83GhJfuODVRO12jyb4bDGYy0Z4wBWk98f1XeKfJ8a9CR/dLpTp8gs
34xPt909mnfPpaB35H2MGdud7rrf/tYXFcx9xPkPAwTl5LB4xwmfLPgpDYaCdk5RCD4zp8SSv9We
xM2AzsKMi0xVYAIso4rGYg6nT/ZE3xU1PIndLEv7QrenHy9DK4bWCMBEVMAg8609sdmci/FHzTl0
y96NyLV20Oo5fT9FFxRurdfFT5/R3IudCHJ64SnG6O3IWAjPAcVe9N1S9PnvPTOzRtTGCJmd4H6Z
NY/mAzqQFNWogr41N7bgcEbvfI1YfooSAlK5lpH2G8O8dqgWml3yEO6ed33d6pGWOtAcN32ly+xs
/r1PSjvVU38ca7Re+xWpuwvEqBzplzHIPllyRD0G9n0QqF0FJ2DvjOdz/NSYHlR89kgpipYZHvCt
5ybEU4Is4fkg1YBbsiCpX6hzSbgf/K6m01NOZvlu3v0veTdCSoGBV7s6iqG7z+YsuT5xjvpkIlig
s0lYZPf+LV6qO+n/4n07F/DiZYPEXJnqe38MnsiPO4Geb+AVgL/gG/Fe4jsXXdbbhOPFJB7j3Gj3
UaVpcacdv7QBoC/kxvNYOTbs9N+VU+alYliqEKtdCqRRwlNA6GoQo7OiB52bmnNv9G6UikvEGPLg
4IkxsLuzDSHFRjRRxz46mPpV3RLC72AAwZkXa8MSGBXkwhrKAsuI7Vyz8SXCxcxYJnMxyTarzS3M
5ihED6eYPaJ8aO6nleYDQMuFkg7BFcj/dpwbzwRaX8ISUpI//y3B7AmTPYecnSlxUHLld4wDfKMj
7KFivwqZIbtQS45nb5D+GSVamMwjqd0lseYRH40nGUE0O7cFcxZqHEbV16zTMz9tmaGkDvfj1oY4
RfcmG5LhbnuSkYyl/RO7pb/8CnDZkrjle1CclWo5Lb8HJ+NYAPSlrNX3R+cYZ58BfSw80qPJDc3c
hqLHUgBHLw26Y/a1Wp8mO9+lneER/M5eedsCljT7LFBoNuveIDILYXDLb95mqaazXVZ4dOsqyEw+
K100JoTGpctFaSb1HLY0eaLfQXX2n6tRO9CJ3g0wVAL8hjKdDY3xFWyjFFdFpct5+bz9wOS4gdSf
3hPJSxNWftDx1C9uk6Xy24Zaf7c1U7p2cK0xEQORdD9xEa26eFEQbsZgMT6t/AMPpcCyPF7k+Ady
WbHh9nuUMeyWRSmJsKRObzTPyouSLh3MdUGqkia+wF/3emPAjLAzafgDErqsmV4p58cEG4oyhM7Q
ms/3iYz0xbvYaalgnrqNh456C9HBB77UUPVVUadrNcgSEXC7LnngBwzZAPZv1itwI/GAexlGfz7v
3KsQVsnbjrtQ7NDzxrfB/89yii3R0NqQi+w7AdYVMEYgRcSp5eh0RiLMpiCtOZ8QkuI0ZHrPfn5s
i9vfi3eIrnTeuBj64KvH8OmkAFtqajKAs3Qjv9udq6O4hjwCyHb3QhPRBK/OAdSxAfcUoiwpKhaN
Dzd5j2Nth8YG7JHdPZG3tRvsiTrmjgyFQ/lnlA7VDfmZfMgDPRE6ZjjMO0Dk8axL56BaQhnz1gGr
fCJMZADbfnk6bg90UjEI6caiV3Dd1h4or5LZPzzakf9gDBAyNdg4pz8f78e34l0Q4EM97OiNJ7eI
AQMoVyQBsuhtXYKZ52RBCuqlaqKZklbJ0SUZoq0VgqHs/E3tNnprjAQlHDt9gwcBdvN00xIkneJY
T7qCwzN65nmDVJv3jdh2h7Fsdi8PU0UxiyUzsR5JqM9sSbEz0hnHy1REV0RYkPuvYEUOHVF2R6Pr
dCuhPWgUvmdLRE79uSwz+whlXezb/JmXDH0IiSB2QrbPvZdcw2t7+kuXGAxryncT8PcwjnKavhsW
Tg4TPLu/jOr7zZJJoq6WL75+msLe4RGGI5dpS2BBdmmZTEFBEz3oxeLfd3Ht9UgkPIGrUoi0S4EH
lLCaWkV+wvxdnwIPXH3c7DuqVu6LIrKyEm25wpek1soOZrl+MARJVdb4+4MIlMM0TwiTSVakK3/R
QtBOFYZnQhvSB4ujf489WdtxSlhcaHeLSJk6oXHDCrzrRu2ykHIld/4wH5MSxGDaRUvw5I8eoz+A
376Gu9PD6W4id8D/PHqQOMotmufZytUnimOIJFQXdAQvaC1/9bkVdS7JxYYcrmclwCV2x/fxo+JT
x+HpTk5JaG5RCJcnNHzYvl31y1XLGM6t0hTapVJWYd0WfyUrRYiUyy4ALto7HWPiXlDpQXODVdUc
Rmb/Eku7h9vPQIFPttFM9GeZUfAA0Bl9ZZ/UvOpLMG/9GNy/D2CBLO5TYC/5xE/SFER8rW0jC121
g470zcfYb9Z+QvXMjxcCDS1qGAkp0naj0Z4DvjxgATffjQ66ab45v3JqlxqDi/4ScYleL+cbdSQy
Xzj0sqFwrvt9ymqHOXmYrBY8NfBSZ2Rohb1YiPJKUx2OPuX39Cew8e6gKvkwGsdX8Yk87Qv68pDK
X/vNSE0WRduMzC5ro+5Bi9GjZULbNRXQmwCp+wv8eAwWtHLtFyFelRHhHQhB1t/yApq6EGAHWlXv
UO4dwjEUv4sqYQMXVztIrLJfYfxkO5deZPb51i5dBVUkZqEZEJSc5Rb+kiX1o/LWEKWZscWp4la7
5Dju9nDBUyDPmNUSPcfuhmFW5ZnJUbimmaPM4xs3QsE8zW9Jid+v0sXaga1R8VWV3Hg//aaX0kYm
cVpTiiUOwVlvF7pDg6i6ZK6zSgBX4oMhlXTG5n6SgPQ430E7+G5O/StXO92Ohaqj/FC2W3fi748H
qxIkTqwtruW+7PM20CE8lVi00UDqgv848d+O1oSHjF4b9RmcJD9nbGFf7oDEfQWusH5+8LyDAf3t
aZ+KHZ9eI5ImrD+aomrnRVngM+adOc8rtwVaA4wP2WjtqnWOwWOaznS3uWnpsm4kA4UEwow8WsoN
u/l0/aux2uZ/RTkNppxiq7QKQ16EMzO5gfsUTU7iseVEJJvv9j2zAUxY8EumUeQI0dZUN4DpSYD9
Qdy8RHWYSBTUXRvUAcehX/ereSPL/tI9Dtsb7dKBGh/EnuRK936eaM+plMc5PkTJN9d7i9Rv/Iwm
j1s9rEIVF1g86MsSu/nBez74dTygQTJfWx6/UBviJnIYSr7Cl5OVruGXR87pnrh297RfgnnwH+gK
HC/oYvdYnwflMWpR1mQiZtvk0ZV9L/Ey0NX0EPnEKiJdE+juaDBvrlpg3f7XJEfJuoC4ynnClgz5
9NDBnCBDcfrNMTwVJdWCwjnPiI/SqEbbWSo/cd0K+wzkENaShpQCQIHiryFZa17QL3B7FbFwegVb
AyXjkgYZvWUHooBKjQpEkQ8WrELl7LDLqdlwA5vQYTSIdgjvGLx678jchT3dKL54QbFDOpgZTgiZ
OKZrrdOFYBoAm+LFPEUdyoo9YBBsyrevEC2gtcfgabl+rr7zIw7cipxabmwJBFOjZbjuP8Fo5w32
93EcUNgBxHnqri0lcGfJqbjg7S3+iv+mARLscM96MGKWKBaAG9Z0FKJm8jz6EPqNM7ojbyeChzBn
Vg4nHiksCOP6c6ryIlc/BDKs+1Vx2fZ3BbJSQRqGgNEIC8ipPmN4+GWe4aU5Sw61ittN6mlD83KG
INBd520iGvgvk8nFODdmXMRcxSqEIe9YZQxlVvrvvq4bHvrLD1A2ZhBnRs8wuQmwG49OF0W4kgcq
Ec6mszCBLAd8UygHkzXkumT4Bw3O8JBzgHaX27u4JtPelaZ/nQ7r5HhX5Ixslw+S7f7Y7fTvPPVu
1cIXsn5akJeWN0UXzA/tK8ohrNHeKpxqVHJZcnEDhPrl+TrCW0+kRboWK+w8Hu2xWgmLK12qXAiz
jKDNKh5KmGr0n7VmWgcavWS8L2A+rO46GgEkBp4hb5u7zH7hKtEh4LJWgZJXR0aCUDzvmPniw8Yf
XLxqq5oW5FyubTzInNWgIVYcSd+nNIglI9urM1/gvS+JbuUq8NYNg1VL6VZgGfoeQWXBNtrdxfw7
UunVgZHu5WUmtzgIvVO2vNREcX7wdgoBfzsJZ2YPs0tVxETSIJpsShrnb/TO6Zsti+RAsZQ3f3Kh
K3D2u6qv2lXCIsnIlCJNrIy0fMZ7O914KPvrcZbOtRWhvVXUgfPIcrANV9JB5LTrlQrcqPH9Qjnw
OnsXKX+sD/lcCnB2wb6UP8kLRg9alwaNAtvKDU+2F9p33fTvppe8yyRxb47zrk8MRlBLDWZun/k9
e2BD/3bAlwRd4g3GghfVPQFCG3VIxaRYydsQ88uk3ba9ho1s/aPNG+zAj8JUyAaFepiChyHsXA1H
KisSxfUMlqRKKe5+Q7pSlhsO+PzWKhFFiWLtuAMpOnR3A1oyZ4MYkeRrZQGFjn7oZS7p7QxkuONI
0q1XNX+gVB1AS05k4h6H2sIK/LGq2RjJeIccX9ZDFaxZXWNuj0pFMA9Pc99vmDXincoadJ73buMZ
up/XKkSEO4EHehRAzpabjyjgC+8mtBM4SfzOgFvmYiWD3ZIpUQNGYNXfjtOE2gVvO+/B8/aKvcQ3
TJE5Sl/H7h1Mezjk0E/rIGnDgKXDwsJtXE9t8Wm1WgHfG2sO4HUxS0fyF6Cz3TN5vp3jRqPJxWpA
SgO/nwFBnX5KJnuXwUAHjN1nrIP+oQgXUWdVNR+LTOrMUNxvDeOeEUbct/bJ6WnWP53Gxr2vEzZZ
Jq0KrtbWQFKI1GyHYneMz/oWMYBD3vfYsVah4ZIvVZFlWLoYuhazygcQh8W+PEw+LxqmqcEaO0Dp
eYbQPWfJGqsg+M7NR+CDIdCxuqMx6SFROxZJTAewL5/bARG2sA8oBKNZDQ/foIdRLnWB/XZdpzXr
NFdoacpMtl1q/FOw/ScodNYhKLdp5KdMwfOn/A38vfpAxEmzc2mUZtzgiI9dJNCXHTTDh6cDt0/r
k95TexihU3/H8RyZnDG5G2OeZVETWPwbqsmpQbxdkrT60kQSyrJBKWp0s8n/OTKBBa9Vc6vjdmAq
gc1ZFa9BkAGx88tGTbfQl8V/EmOw2nylzs2YuGBEP00mezTRI0p3wi6qDnDigEfM+6kmli6qL4tP
kZ5/1wywxtum8p7G5CAQNHR6tKuNx76IJzECGveXTG6wCWUVWsqNvsSacERbtiao891CfwGqLCnq
Y2XQ3zdlQTJaC4XI3Pl5RTQn5UGcVLwAZaXqCFREjW8gQlx6L4ToYP5FK3By1PHQZGMWDG7UUtZv
9UkB8mgIIxiD1F5sWG7GBNYvjNPDVDU6SQVDArRi6ub2X4sZzghknuvSrGewYbhYOLcG+Yu/myC7
2REIhd6aH+Glm/5NXFb1BrD77Da980WwRlCwo7URLKM/R62YQvIif6A42Q+5URIJ0q6TwFNeiAUI
ixpy9Q/D27q362ExY6CkT1LWe4a3YSFpjEd+SCfcJ7OMHUVF8qtse6hfhNv8fu99X88Td067o/P1
0S5SLN1xPoUBJxEhcm1z36fb82JI59VL0aTlnLeKUQWQSPAf+bCSjfnxT8ePYRsRvxPtP8LjMl8X
lYlqaG6AL3RxQWVgdYtBiWS82rHHtlDqbXs+2zwybGtD48i0xOk/TlJ0ycAMYyJojQGVQCoADCuS
5BY3R4O851gPdVcwBqHKR/CoEZ4shmwUzdc5VJbylCmOl/xt5UsxvB8uGjkOwotkLNwXgVkQYX2g
y6iYCUOElV9OsGV3/+YcreZhPfQW1bGDs5lwkndRQobfUyjw5OivGlmiv9Ot4J6A1EksAFixbJz9
idgi4QIdaQ2DXi5/Xz5uB9BkhR/8o8B82M+vQqX+9sCXryjtjeFSLL2Sc9hmTL33jb0uCnmWjnmO
8u3yuv6u+mjU7uUN1JreTPJyLXzGPQ7HO8m7CXjYtwqxr0+2iaezp+smZUNDhtyd7D8VFGS3qa0z
ut4tnRrUgLe6RIJ4lqZLeBCgy1la2pwlYITvesCGpI1jQwd0GMMEw+KsQj572s7lgAFrmuy9Slr3
X1b3KhIyOpuuO7JzBwK89+FFIu4Y2ZwdWEuI6YeEQfNZ3s2GtexgEVEJW4fNyL5Y9+KWFqcIzGov
DuqMUccTaycK48gW0uR6H5t4ynHT3rdxHV0gfQlhmtge0yzyUn7cB3XtaGPQoF0EFtNHzy04mS8g
DgXiWlu3WE1ATJwy55P1jJ3PD8qzFueIIGTKsU4NlkBHDXfHf8fNIxNnBHCFPfIQWQIwuWI9KC/Y
/79sHZITpfCTQg/wnJl1dMjCTH1VvqKs7+rEa14LR3Byc8615mRigx8MfTCYEt2tWAIzB7v7XWTj
T0+0jCrNhYYcTxEERyB3ZbueuPWX9r3JFQ6gVGJAEzJPMIKxrwg+clnpTQ173Jhd1Xj0LRE0VskX
wWcTbUoqmXLJFa/3JqQDwzB0cYwWWdidDi6dzHaXYFNXFBjKkBlJjBCAOqV8eBVoOuleW45fuKn+
y6WkxNkfDwqoQcYD9wHh8xF5B95i7iEBD9A9+Ue3aUlYjAnvufiJFRQhInGR9PdC/I/muYQBxfA+
fI1UdK6/HRefiS+FJIf81UGLNTurptqMeh22WRqIlytXQocD6r8KHH/Y90jrOF1XL6OfdDdC7Jef
0LV2bjK0Le+UhkDGdKPurMCWJUppqCk7cSzTl4BGFDRE5JC9OMMQe9PWEPEwaVWkf1Jq/t4JH/zN
qmVcXx5BBwyql8k+T4SoqpRb8UgAfina+q57ZWeJh0dArdTiqy2giNMS7ylYL89q61u5Dy3kwiXS
utw8Du0uKb8h8XJw0T3WTQ0FmDvsWrKk191ru9vLhQswDSzB9rUvgYLFSXMRW9n7Gd4V0QgduSrK
eJqb1Qqsr7AI/y5LsOLQww5o2hvHIopUuMmSbL4dGyCWX133jm7s5j4lrJyt0Z17e8lD4gWYujrX
mNdidl9yIWmPZcWgm6gP2yj1WxDUF2XkaMySzBIr7FOPpHLKYA4CCdwVTWhHf07HM1JBSJDa8Mxp
/Fd8pp2zUzRsc3hAZM59l9tsffABzX6gdrIFA83K4piYHwNnHGdBd/igDTCCBJY6H4V/Wqrk9Krs
kbxr7hrqTn+kWgRQ2/w3YQoUFc2W/1myfLnIce5F8CCqE36hWCWS+1HgZeFyLtjj1lj2r5quBVh6
9JYVUQAuf6VEjwrqVBg7WciJqdNlgspjdDsv2wprOygURHgm1crXhZcv5/JvHywUv2i0wm6BmnXc
yoPCFUKRij2y8CX2EyUKyy/DbFW6bF5yEu9lpCap9MRLngMnHN/zgAtovpnlL81dBrGprBI+bJRV
MgVuf1yj5Bf3VSgT95O8iuYDcETmvqJe5DGaELcnkVDeI7v6msYN4t3DK3LZtzIyRJYsjR5eDARJ
4G1hr05rgkgy6Sznn2mTPw/lN2Si9/Aons7W+nN1cfCXlyzGXW+604go+qmWMZ5Js+EOvBzwiZ3S
uThTkdf6ig7Dy1iFm0hlygKxdFX5+pYMyaDmQOqQYBkJoviPJcpSaaRvOKXx7erPQd7Bq/MqNmei
tFBRvxhWq+MLAE7VX3+Q7smwq3wegq6qq321Sbr+vyE2Pt4UfkdzD3akdoH//uMJcQnuPaZNQ4LJ
MaibxGU4jr7JkwpCLTgjtyLhNCoZSAVrSLiuCLpFerqeEbfRnzZhLC5bdGGWv/dkJ0LG9SfV+mE1
H3ODaYgSW+O3/+U9O08P/T916OyTUUmeL8ao36x4krOSI/fw8AtAr75oHCuIBGi0a+Hqz5zVcmxY
+ea/UqGl35ZYzjLCPpRpcEthviwUdPKtQdKzDjX0ghgss2EYuPw+qTuXHACwzjW6oNoeVF0cD1yH
2+5Wn8XZiqGP4jP9Sa3RqWu2MAXgQWjBLTg5z6rgDcWczwtYw2QvjExl/WaT6Ho7yzJCSRV2H1Im
kQjHJSIDH4h4QXQmWNFAUjx7ptDbYfFZCdi31SnPbozhhqFTjtCwL4jncCxSUgsJxSrigysSzvaf
Ey1uldjtgDebfZm0E8Q6XNuH75E2hc6Uu4kxkZGba8n+VPm4vfougR63SZrFUIrIXHhcJAoi6vEN
30KW2oXrsMbP43Sn2gdVKUDzRbMdlnLWBqUNYgE2MtKu/PISjR5Vth1abrFP7wgEvyJ2gnanoIj2
4tJQQ3s4scFl7CTMFEhu2HA/KqrgKoZmgSklXCyQekeLHZxogzxiZBMoBakPFUVjZcKnv5QzdXBk
9jEdutSK8plmTRljOsGrsOBp/54hJedMfcBCajsCpGvIwVSs9at2o962PjbtyznZ/BKg20vxzQmz
4sme8ZMR5Sctt0cOBEebK4cZYk92Ln5HJ2xrhCS5racHlJy/emN+JeiRNQcMyTbHk3qJAR+Vk6vp
0HvLG8mPbJT6gRje3gJOIL7nid4C7HZoGgUDR2sY9tAF0pwNnlGtpfJZzhOScnerfEsUjXhbcMgJ
YcfkEjZzNdADE01QVgm+by5ABCNfraaPmWGL1bllxTSEcLJm0iRz8BWCN4EFxSyAlqI/jG6+TuSu
MYyfUTzMTNOTG2h6zsiapH+vKF/I7TMtV7+VMfyro+EjshfWLe6iHt9PG8hVHpSM7yrLiPOIcXRV
shqN8UgTsfOIyYl5UxbUK3ko45ITt+xnL3Cp/hFHl6MnkjKWshotJ5V9uI+IgkeZaKZDUxkWI45G
Nxm4eE96hw72UXNjNXnD16pCyrbYjUdZ5CuhaTpAfM+QmRhFzdBSiov/Jj/uLQwzDNqoauY+45z5
XpDz0Hcf/oO238A+/slLpyvIK1u+Z8L7gTosrUoO922NSckJj06Skfb9cV0qSXpPkr+RdQifsKqg
TbVmdftSxz4erqnfSYb60czyMruimly7bQn+IU/J0maItySo+jpe2k3F5gTkB39w0suBqUcTx/Kg
uxl2f/DTR+cnCAdquW2VWE5XG+Ypf93WxjdRVpOX1V/05MYtRxRuWxxi1UaB+Hbe+QNzakcNBtRb
LlGifi5cOhIsUiYHdDzlfyzJ1lD3jdEHd1ZNxNYiqea+TH5r4kmo9WfsH562rvAuIh5stSbTy+00
vBU2x63l1rvbh0pmzZoq/SiOhn16JUWjEvjCdfUfvvXXhLTCZMyMtk6zOl1UwxV+rkVogR6X3Vs8
84A2b5XGwVrnRaL8PSOQewM+f/ycMLrJmr45bNPXqU2xnwdFHE9ywlLawHi5SwKcnWmJzQnJE8CK
f55W9ky4qSztce54GPzyWEUUX3eL7DDIZid4tqBrbn5Efkdpvje7PvE9byMfECXZWTl7T7lLvta/
zSChQ4AS/9bo8cX7ugXk4RVuaD0p1JiYHmBvDjVAbKAdKGkfT2wwH5cpNQK+HAP2fSdj7MuttmZy
PHNsBqUkixnrzcdHl472LMI8SftK3f+of2kW110aS47NNOxdmSHKC3vEUxw0N++NgaKt9w+nJnYK
3H2AXteWqw7QMA1IlMF5qkgKTZCBVREDB2cE9vrXP0mVdTUiY0sASprxq+YCeZEaPpYhLFOZl2/4
S71WjNOWSfSoW/QpZIkcK0mkU/D5YgqynnZJ4o/0Aew2q6nTzBKt3tnGt4Vkpptq6mf2uk5fenpH
Pz+oc5oNVFXNXqGnFna47dIoqt7kSuV4VQ9ACO806y/mKX5O6mj+ipxKzSnN9ahydjRDqXWGBDkz
LT5vVDYOYzMiUN0joauBMhxyaguv1jZgnkgl73vMUlkMjadPviGwnLY/H++rIfduZfXtxfir7rwo
I7MYYdTKzE4rQ82hglvZIwcnps6FnuWigFb1rRIR6PsfnL584vSPUiGAzOfsIKVc0LAkmfepdrrO
pXvAhWl632t0UjCoRtJ+gF73ce1L7oZyBY0MDHKxIQ7opAI/v9ZQehYeJWrwXDHtLzK6ZsIBe3Uo
ElQaX4yTEpKroTrMnt8BEjuxI2NB1cyV6v2cyH7QXzSDJKTIBEdaaqXAN9PB/bTApSgno/8Iuxfp
hpMWBU2MHSZrL9y39+RNBnE6O+n/bqt/ExxHaAkI+oUZBqQxxG2t7uBNC/jfXsU9SYHaNT4jE9Bb
Qm6XpeLJvnMoM8FK9lXitHe1iHM2g8pHSkXwZ9kPG8+RhhS45T4Cnv9nRG2A2ZXttQMHOpexP08U
Djgg9S/xo+nXpTebo+WB87/mU1xnAGjSDeMGAM4TssE1wzf4HLCgs5TcQSGrdu5tYY1K/L7hYB4Y
NiLWPWWFusgzTM8qoFuF8NJUJCBsbaRoRpcekn4+7MhSZew0nlzM7SDjCCCub77ThkTLP0yKSFuO
FZzdxDq+jNL/qov0wbiInuPN7CELQ/yPIk4mgpuafPz1WSgRLxS7SGpFCvYTf1uiKZV50XD+SU7F
ucyBiZpaWCyrZTLJWJzc5nI53g0wOhPycR+sSmxRlvQDWmdx/U3nkRTiA28HuK4HzDR043D3SkGB
e+lb10wVNjHea462w2tgC3X8HYEsNdiWyqmPsCRaWfcw5+gqwdXS4DkhQkYzVo8F0Eptlhh/jHIy
WGkrRVAaN26s09YfI4ip1jhhMQnwaHj9iA6TsFsgNRJ5NL1efEuUHJh3ixs7EVrxy3wgYXlE0TcG
uEuWWsVJEmp1M//dh+Xb5gk7GB69QXl4+5w4mAdjTuDBLy/pSSS9/0JobDk+BnvqKVZhBMiJlpMZ
Ku/0zJ5aqSAFqTh85l7VfCZv2eHJJhCcnj0+rK8fTP0u+yOLAIhmqnpcyRS+SFGU/0cSsfrNdSLZ
DX9Sipc4wHajtv84GJJTl0eSNoFz0tZ7H0ZNpjzsYNKU4X4vPaMfSXCYBfvZkiDTGQMWuk/dQvt8
5EOJ0oGX3ei9NUaKuR9igmEEr1y0hidD6aBjwjsaodfGaLxx91neQn/ubVVsvW1moRFteOc/Kk5w
snSlEnBwLppJbUawrWhW93+8jvZZJI3O1jGIb93cTELgpTE9JOsT0bQiI+uY5xMvOgG2yb/4SrOP
PVo3es1pshWMiLzcaizLBoIB+udxCNtfoQafmGLYlgemiNorSJH0T68WXLTW3+gmA9GNdq6xoHhr
5PTn6dKBvJq1njJrRN7stNMgw6oWyHVAeTXMu8BpYPBU3J4f2eeYZvPtkGEJMZoJlALIYIzS5+yU
jMOXkDVyHcBaSJXHIqFyeAut5KEYeH+zAuHIKZmv9BwmbqSGwnFjwj46WfkmIupe1NRRx0ByYBTa
w8aw/smymz4sDc+y57EsyWz3EfAzwngjPvh8bGGZyEWRxYcoJ2EZCnRLFgA1KgB7jTBBLE5trFfE
+FtcWf+cyq2KOm28/iLnfBhKT3crUmpj0koN/Ux8ZqEj+Vyp89np3bC454RdWRj69wlfXQLx941c
3j4MSqUkr8gJ9iBo+v/ZZ1LeIyI99/yX5nY+mAnaNQ5kPFCI/1y4hIH5C204+j9IhAOOotD1KrGL
E0zha1JQna7OwJl6hvP4yTab/V79szmPX+BKBT2/wE/mCwljdrvLTG1WYQHK8f1fdiB10AsNtVmb
LIf4ibEtKE7PHQSpSIWO2RF8ZwBVp04vjFT+TYh+qs1o5tG4s7cVHaxgU0W3M+pV6a8uvZZhO0sK
WDlzUgaREpzpCfcLUJ+1E29PrVZhxoeAm2h08XTual1W+bmu7MDs5OyakacxhdmEW/yCbDZefyZd
YwK+HcJW8GYkfkz5KCkL7DpcbRvM8pbosccHpdZpLKajcTNs38XU7u+dq+cAK79uQh9MeS1NU36V
zGyK6RGUsmFsqgWuQE388XzGQ9UFOiOmpYNF0JNiaIWWV0h6woV3MPvh02YzHdo0wVpA+qjYuIBD
uAUT8r2F7wgPhXIHsVQDe3loDc9NGoJPg5x9YjHY60pByzuFitlF+ihXEYbPPnZqrheFtf4ZcFWx
MSo6MZM6Vwn5e/XHfyFFibjFn7DxCYBBGekC8RTVFDvx2ay1TubWp7GlzWJnUaVtX+Aaf/4uZHq6
QFbYb3+1jqR5MBFPwBJ3AL2D1ZMEkN+sBOBArF9/wwpCbZCwRtS9QsYLjp8elafPYFt6cz8lwXS8
TlsmdyO+1htfY4JSQCIzT+RQMGVmFrjCd6LmaZaxQAxjmqvBZpUnSFZ9k3Fc8GbPRJaocwqNsWSY
zi2V992qJ5oLtA9BGnURgjD8CtSHeqKTz9mrHyaPspaNcuT3J+jDAsDJQYnEF03V1B2ja85A/b5A
iBttTdbs+Z0z7ELIPO348Z3uaBveocoWY9Cxmugfgu2O3ggRHaAgFo3nv0sgogGMqaGa1iF2/9Bq
LYTfZNu5Okf6qAwcUUp5JFGWEj/IWeZYE0UxDNRPW35eZUl4chk5qA+HCBnGHsaEciBQDLphrmmZ
CF678O5TgKrqGyJNzMOkYPX5Gwv9x4TE9CTvBwkaYQdYq3xdU5J6sv8S6ghBT2A6OoO+zOObe/4K
doxxHyon/7bsO8DXicZqt/cisSL104oZJuU9EMsVBn3FDbqDHHobaCc0PSSASo56nKZ4xbwX6FhU
M2v4Jthdsz6ny0RrJQDyj34vSfvgXGayDj/HdN7uJSn+uRMFGM73jzXl53yIu0ueRy3xDW6byD53
cnwc4PU2o/8NnFYC9ivObdHicjxLM3+cjnbOVypLMm6tLvcmRFRZgh/EOpSYAlWALUg2DNGGHgQq
+dh3W3b7RaQ7V88T6TjquWtRD7nYGAImbh+z3SLHTs9Lb7ZHKqCbw2H5C3qDcC2UWijvPuGYkaSq
Ze5sdVK/x7JHD9y7b8gXXt3K0qxAcGHRzng2VIYaN+Mer1t3TiYfZtxYaBIOva18MBRP9Yh8L0Mt
9PHDkI874eUukMYx8Y691GNrU7ybwiR/xJZQJYmPbg8297jkNRug3oGB+ukIYojNSW0EFNK0Q+so
rgI9UKYC3ES5QrByXfMH8UAEQmdF4kCaT+P+iGu2rKJS8Lk0XGh6KwM80aqOZxtAyh+JXQpU9na8
CeW0mFOJb/f/ALnVsqeZrJBSdrYfVZyYUWPVeHhnCte9On4sRiPxxk+J/iDbkSunI9Td8PQoWkoO
dbLScHxlhyDIQ3LTuXNHb7LyWIiUvVfZ9ed8NnQtUy863k3+hZ6uO4zchRm8exsvvFgzPjXZqAty
/Sf/ky5nWTAciKUzwWE9kGemrrZaDoqZ4SdA8GPwiFkhlRCoAYToYylQ0iiu3NPa46NlwJRZCZhG
KRfWNMWUmX6zNpmXrKc2Xug8kPNUL+tGRVdL9c9b01pObys5kgP4WG7bOFFobYkOGPB4hFkeD5MU
9Daz+b3LQW0uYKk92riskDY6leRMZ1Z8T2iaRMYmC4d2Yuge2ARzWFV9bJve8C3cuau3BM5gEA4p
H/uKMouzpsrA53oITdcjg/t+//Wk35eAseklAKvP2YHpq3MdU9+gZsDsZyye7hDtqgr3uLqdOXl6
HbTZ//VxtytVsL9Ld1ETTL9kTCnuOSMA5htETBdhsX1MzPqpEn7NrlwT4khQBfkORoci0ZSMhbQ+
ohHCUhSoUblge6c9I774SdUZnBlJNjzm3AOxqPK61cq1ISWckkBq6NvxGS6Ls23VgV2t4eCXex0j
cAjK/HNqANHV/NtZu6PAPQajBew91O9u9kv3QEz6QFA84wyN+l+nwfl1LnkAj7v3ycWjCWMdaPYX
FxHzjMjQdsMS3XpcujmSuzh01QEcwp+0qbSJNtjM9dpGTIvZD+wXZXDMih5BnGzD/Li8Ncib5yDz
qayGbHcLSrKfXrOFMafWmEegw64N2ucRZLRUmI5lNaAvf53EgQINze9KvB4J0By8GPKVipXvHVCL
miQqKd/yBQOztk2sz6ApprK9xUw4KMnsGb0062GoLWCnwVOKPVZVte5AA1JIwz9WkxnQZzJWtS1X
uw71fkaf8MeMQ96cdzRF5yUKOEVUgjtNmvkK+kt2b0UIJxBa1rSl3kG39lTuMlIqerS2Eppcnynb
A4GEzpp/RM4073acJ42iJrAyPCfnwCSxCTu64kgNuGjG3b0QBlSsWdBMDoev5SFRg4Fi7fpSZ1tJ
ITr+e+g5r80Ff3Hzs0NJHzFsxsO7LNcc+yTjBaUuesVXN7FIPGW+VwQvlabZBaviMeQtkfskK34y
rjiPa+HxQ3+ivlcFwlkfxPgID9acaS61Xr29ErlqXu5oNBRPlrfCdiHen6wX0auAANM/4GGOgKSL
reOqUAUaU05PeDtDjmoEbVvLtA/6Esvx232WgBTq8TyrUzI/x4SfJzXj6rKfwcGtrJWxU2jBc63o
utQr0jfN5wxKuR3J/ff1MPweP9KX8Sgd/7fXVPYDH+HGql63laY3dyEUfwUs3hYkEZv8UeZnHWpr
+NkHO9UVV1cYlzXw41nV6jGC66Ipd3krqDDxSxH5LP7DwK7u5iNivwqmIKYboIFExvWBmC9maji5
Y5vjjuvH0rqOi5/hBnDZ0bV5+OuFj8M2iVP4Cp6rF1pvTJ5FtV05H8LxhzRXkRWkRcyeRrV4X5ol
9gckrIFzav47Fv9Xyo+Y617i7ZchL18jsM1IdIUiCzMcbP7375hsZIxGNEd+89/Fg1LbQMIDf/MI
QWQK1NS7wFSX9kv5vXmTMGstTjdJmPG0TKf4lvUPkC3vxEEf/MeeDYJIFQE+SaQ8Qiog+NPPgwQi
fxTsoVpSw5lM5CQwY1/0D4pwJrkA6/VZ0VMizYMs3mTKZILde5EfbW0vaIe++X1y/LEgrxQZ69Qj
POcMn4t+lCI4Twm6qyNyJCOnyCeXscg+H2/KCn4CPRzJyKAc8l+J4XM93n7JyyJVQfs/WUi/1RLx
OAVTvtGS3kgK39xoL9hPi5iMpWf+czKAESB2RsAMuMD+l+4QdwUmIhvqZsQp+QuHbg8sAZJR6kAI
kOKxDRmDc9D+TajabV4aGDZDfwyggKx5FVoXDGsgDgks/jbb5vZZw5ZxZCZLWntZ+Aqa6qOXEcNw
IieY0sA8zPA/h/8BmIFuiKL2vLJN9QcBIgkrBX8VUSgYC922ujl1yxSSpLMTZa/KWka7HvmTANHo
CLNYo6eucFyX4wpeg+gKS1qjfVnDyz2hEPh4HYJ6vXbqg0sJxpokESZUFG8FI3lm+nipbLTZBuEq
YejvDoGeNjRTGPAW1rJTOUtuYQbu0EX+mtd5p6JB7rBRUwN8T3NglRayrjBU9anicYbI2xkbjZYk
RT8TK8hylqpvOBJQvEnxSLR5V/secT2Vgq3nYKFa/nf8HMPs0v/Gt/8hgNgXMbW/Ym9706IfMHIQ
7f5Lriqm+nxRVq7itF17VKirLRJzAdcZ+TudBrldubrbf+gWpzXvesgCM19In085231V2RLxvJOk
7GmUk7cp+cpLsk5qShJ1rMqrnd3hcDcCZcUGYEqJSTnj3+DWesJPDAekuWxOz8TDObevwKGi2Mn3
MzHw0TsWsMZDQErIjnLtFxx+BcNm/2ybhyxIU8zHEPNeUheEgRfBHW19lDfui/4wuF6tvbz6/6cm
P5Ee2CE3Wa6s47vDtlWjV0b+J5gBTGLXxfqxDO963XRVavnHCVozKrFuxAjUCWPhWOQnYVqDOTyr
S9f1F7YSqmh3NdX32kUhJRV82XcwmdD40EYAp+E2FDK5j+54tTtLfb72mU9hHnhOkTLQhKNH0pna
202hdTkbS+fG7aiptHo3y/OysVsTb6Ry5AwdbtEbJe55q/aYD60iAUQCecG0SPZmeN82mbkVF16d
DweO/ln85MVZ73pJauSHaE/l9FwhSPGru6i/2yJLiWu5iPNwaxonzOiAoMnnpnVt2bv+fLyXyKp2
TKdg72BZj81HPUvTe5zfk2LqZhcZQ2dekoFy6cJXmvOIV2jNswazQuwJF/Cug5Ic0NCXj7pMEjX0
mv6Ij0K69QXJ3IubtEBqd9+KL0H/B2GHt24uLCR3Ger+j1cRF+D9EFNUxbqIJX0e6RHHBa+1Plkg
iFnzmvnicJdDDDfS6nlfV/53Uv9jqPrU8WfNQG1IF/CR6dLb5+6Uv+vEsLlIAPIdN/vPf2UMMD7N
Nlh0VxWRhxXfbDmPkYSimfOFvVuY8qDtYiEzhYN62Izzj9VM8TceFB97I00r79w7xR045HjekV8I
h0vQuXRx3D9AxelnNqfpASJclIelFC17yKqm3Nnmf0c9q3VKNg2h3C5HPj0hf2aonY2ZKnfExdX4
2PGCLYYc6YvevbObdt6XN/DhdOfq5ZJ1c0//Ebhdq8qrER1SNl8p9HMez+G4IG0+s0saagZeh0Px
/fOLaLqlfAn9JXX3y+G8mHG9NM8Dtl8joYI646VqMzSPXTJTKe/oJqk+cv0HoTOUGOTcPzXfKEma
zDiB9xoxg/4TEEA4Ckk9u2ZkQV43/CzFHEy9K/GziqrbJzO7ynaM/of128e1lFEap73hJ3rxvxlV
058dFhWpmbr1ZdNe4asFlWk/rlH8ZMOSTXLgUta22IV7NNIEfBYhprC4l54vstY7FieTbvD0izNR
OGmHnenqX6YfiJDNqtxoeOgD9xcyQLuPkeNrWjEWVjb0+v4PJt2RsI7+WW6iHDGrhoyEMZxoaXa9
DK3f13sGr01d2DHPgItVLZfSHHRNHFe5u0vuLoTiVDGCls32rsZePAFHAApcNmnSopWHARJq+PC/
BozRClK9gDdE5KQeKRvXLLt6Y3BHfhTHtJoU8PmbjlhSGK99yxouLOVYttBwZ2z8d4GIoIR1szYA
o+f64lFY96IU5ERDjBJN9I0eDGKiRXg/309gvq8hoMqKaIdakczUWqsGOMZCGjs6//NAw3MUA3Xe
Ws3/m18RevyJ8WjNuijzkQ71yWI6groruMZC9Qz0uoJPXTstcdvRC7AWxHEEUI/hnR9U9jskEU5r
MjZiE3KuhaGrjTH+762BVbWoGbuDcPo6lX4razFauQDv/piwk7ifctXvFpntVMUUfpLQlGN3U90Z
IR8yUJz+MtZELRSGB3wvOd18+vXpeqTiWDqwH7nrRgKVXyJRnefqwzaKsxFVbSVpg/wtnhTv0vs/
FCfTHWBH0Ru23l39LIdEAqBGPPtP5j4JcrMT2vQ5BH8sxjH15e5Gv+G8/mOCHl9ObLuhYZxAXyvo
uKe/8JuUf2AdJmbJWTgttLyDo/9RSpcbvW10CKrSYCUs7r0BvHzqfY5psuyb7F5hTigAyvWT1x/V
QS4kA6HkLSgjvwsaFRZiOUlbpnuiRwuFPJPoXj4d8hMwdZMYIU0QrNQMPB2ldYK8pStDFEZJDugx
4IfalJmthjAQO8zUVDPykN8Tjc++VVuTYbfKd8uEtvxp6ST+bxdtibOjHwZQF1eBygUBmOJgHcYv
Svp057DTcXp0eWLMIZlcJsfyocwvh8lRkxQzUbQYNkNUj+hpX6ibz9vYy2TEYgtXyR9gUEkI5dgS
pVQ2keznRLlW3xrtbYpdx7lBautNiHCOYPF0J+y6S+UNkLriisrdhnjaWcYlouXXOk5Uh63FVEjc
dgA7tRSMGkVsJIyfWVd4vYPd0fyeLOJdpC8Bqqne00tWsLFvPB8Qjp5YCVNsRfP/ECwfrHkwMdlm
5j8MbnyfbTGFG+TJvmRs3QKXaDM2mupesoqRvCPr/0Cv+TE++wd6cNAnHsazuPj+1yTNSFiM5ec3
XqR/Mu6BzcNLHx8KmhC1tp7Np0huTjbg7txMdWXFF8tDqWyqnY4mejrHK+gOhSMy9lPlS6iOf+FB
ZHHw1HixHt/OLnRAH9k06ZnDqb6knI9m45tH/L+5/M88E91N0hqlrGyhv5uLzRyjuByijOQUdhgQ
/MY5kIcAYUk0qX78WlMLzxbqdhJEdOpuNSjDg7cCvKG+eDNidKWw2RxmTUVPhnQcTwrQWhliWX7W
tqYZazzQaaq3qJ7SCdV8YnHlqrJHvyvyF4pMOT0o58gStywtiH1xenjAV9ilCYltTbZpR+qLmnNF
LPS+UEcqQNsoeSfW2b0njhUhHCk4XMjLkPOZn8xaonAlgZqQsb4ahmsAayHVyKvnIMjvI47tRqkd
S7MVX6YWgCkAc5w9UjPLmQQOm00WDEUK/pnUDywBAbK+ib4yB49N+SCD40gzd4czkMqea1Ar+P0K
oBGBDkbqdjopsrU8QYWpUgi/I+AG621gel3Ry8pJVKHCbXXdodmFmXgPpideg/4oCCawL0U4Hgzk
Lm36MgjXRcZKkjoIp0h9uXTRzEZ2kvQrNA56qSFEZcMZTjSI15ZuTISE5VshcEG/gqG87K1h//q9
sAmGh4X7jG3jIO+eo8DfK+zhqdL+mRXl3+qInmiLZcHfCMJsgadFMAp4WkzgUeo3GW2rk9QQaQuu
P9HVtrW/KVej98Puip8mDO+a2EnY4nxzuLsZ3vYGIh0Ho3I5BBJo4K6MgYDMcO4GOLZ+7v+5qSPx
+b8o7uwZyPNFNbDtiqPDqF1TkvNvbNTHNJK1mfip8yf38ssEuVcV0jxWpn0g0UJGf0Ybpwtf+KeX
rzsxofC1hJ8CT/9e3jAo9TswtrNNfWukVOTEDKsrvBeJ5J6HvvZPryoedbqstqwgKssiM2mewVXG
aFzyhHcEiKziFWbXEtaJvFv3aSDi6ltvDIUcgp3T0JLAouTq0Jx0GqkjTYgba/m9oc/Q7cAfvAPt
UCfcOBUnw05P2kaus5LtFlJCrSHUOKnKXBmZgSqcpna7cIyDuFLBx/yzy0o7EadwSS0qWfIXwjqR
N0Q1T+9An1SZbEo2q9CS2w667UxOkURJqys4L0tz4Vq+zeIoBrSNnNneJ4UbJ5gfrVJThEK/9NyJ
TX8a84PgZcrx4Ac+L4k7vJU8YpD1juaYNRxCSepNIzRC6YJraCWr/7DUqZuMvTS6BRZX0krhN33z
GfqG1Rzj7+QOEZ9qPhjeJ1ibhW012jYViFdyBSWXbp2zysC6cqwzWIy6xkIM4/Alwpv9uGLVR7cZ
pHt83+I5LGpAb+Gts3/VL/Gf+QrZixRlQ315KTfx5s3Es/MEEkbcik3CBpiR6DjvRZBWokbdHdE1
v7gJfbDJvq2T/9kGGC2cvGD8Gzlcb1XwcV4skw74kq36Iml/LX+XGzaR4BqnUlfQkLq37IdHaxDb
1beQF3h1sT/gDfyeonaVe7OOICnfcLsfB0n5eJi1ZHfW20SquVG+zdbGVuZTr59rIaPlNlp6m4RK
tyLUElK5YDk2bgDetYlg8nu/WBu+w4BIwer8WIPHUafPFM4l6LgsEYOBN1QXfuK3pEcQa+HfuW87
JK2eCO81t/VjLFAxbY7o0re/xDrg4tDWSaR2xa4ErnMgb1YG9T7DirOtNZtWPJir8zknwwBUhld1
4/xltfK0SZbOIpepmGo+gaeG+gaz2kGm91VvMyFH7oojMAdHN96BjJB3Bv4svuYgTcDHGmKThqJc
UxwD3JDqpgC600cZJ7Glas0kU4W8Sl63d5wyjud/OQd88nHBxcqyaPoo2VUhDKEd2VyibVK8JkSD
K7lsvSNkLZUzlUWcqinn34BWAByKU8Yg98lCFhhmO0lEaJFwZt8GDPtb65udnIrLXQyp+r6Q7E73
QgsI/81jK9UFsbC9pFbXASc9Jfxo0gg2cKIdRwDVUamIuQPbVeJV4VgB+6ADNAHPbGGc2XjFiHNf
gcdlzKJIKngHEz122yR5snPAU7YLZaw8MB3r9GYBXAPmtCzWjHKBvpCza2G4wr+t8hnmOspGvF9t
9IE00rI6kHRY8t2DdjLFx1Y5YIgTk62se3K++uxAjBNla18jyt/Sq6uB6xSyRXEJGnGTHyaWZtRg
6MW5mNNIHqtMk4C6zOQUmXL5n0UtyXEtq13mv21abZsUuLx/OF0cqeORzrY1wbAbSzCwmXcwP5m6
WCquE++yndEw3Ce2bH0DxY3t0h2qObMui7990MbqcN5IrmjnYQLsl0US00qeTS9nk1JQ/jtMCyz5
NIxP6fA3yEtn+KPLmAiiAwiWZ8UQKRF2bF7T1ocffzVW1FwjAdohLI840ntbrQN7F13ri75zung3
Kt5ucGmBDnS87SadIvyOBLNT1eZHkjjivVNFjfPOAFLS+LgroiNMilTeqK8R+oloBPMtT7vHv0Ix
0Up3g8AWz/HlhVsvGWfALnsPnKHm4/sG+fg0PEA9U/0aN45d1/Su9qOZ535KuylXf7MctqPYYa4q
ivWJpsfyAgmzTPhxBQz/wJ6nQIhaoM1M84KF7KJcvheo15w20Fkcd6QW+RdFCK2R9CBT6uCWNeTf
9zXm+Jh9HccMsaM7A+ZI1kf0DOsnBxJn+SrjgYMF2xW8lEhAKIIHr5f/qoVIOmUI39ISSb9pG4FO
8QYcPfR8WfwAqDo6wq3DN4qlVq5dSk2rYes92acL2rt+Fg3BsXcrTQYwlDWnsN3CIgmjBATs72rD
UWp0d37N1Eqwqph2VKf1lhRIqawAgan0Cpr6+HP4h6RFPLbov0pKqaN25WTnVRb4NwDTK48M46yo
QrFS+j90bd8ve9mULa+zA0rkHTzxizGh5UdRCL69feTVHcm6aAUPnfRXly1ypkyB2NoEMrKi6Vrq
sYV2G5kS096hZkCttHyVeQXbtJTIGPR7ouaWpncyk9gE8FxjPvymllVEeerTUqsTxjbzHCtHSA4R
TIs9Q58LehlydyazPhI2xIPSUVDUPgw4b2hxOLI/4KSMZWBPb3y3DrGVommuZ21WzAKq69g1pefE
IGIFe892CfnjOwc6kVNPlkdtWJ9bOBiZSBRHt58tPdHDiElJ9zB4HBV8b94UCrOCVxNK65K1Y0eu
AG6IkF6fd2+J2356OaBN0USNVzwer6vNuX5mHKdpo7G/Z23x/WpcEn/quV4Gghufuv1Sv5AvJjr4
/Bg0tg74hUc2koT/KhUKYPpFLyOG0e4yG9tSDH8kfvOiWpKVycrrtIRVEc/PfGMJWoDFWh/jJ/xT
0MCOuBVS2891NYY8Ya4ji1IM4aO9HFuvbNvLN+hD6SQ0yjF9uduWSuu082m/4BHzX62TK099XJrT
mmBkcVwCg6RZT5NLLA9ovQH3yt6C69quoL82quu4meK9ZF2whYcrKbBK4oSdZ4JurWNy8sLkSOFp
7zOidr5xRcYB7ul5b1e53+6jft4edk7trxEH832sbvTisydz+PvKCO9h1tmjKG1u9gU+2bGLvF2J
xYl3PximueGEMkPGZNquD+Toy6/xhga+FpFtK6D0ra2Ie2d1D7X1WXlRxvR9flfXnTIbKxMufsKO
HX8jFRYY5NSpDX98H3HDH/ck2OK84Tee8hi2jmOPhDcq7hPXABAWdbUv6MhFrgrbzBZyulFOwPr+
5pfticDiRgGrHrm6hJn22eVWCO6cSc2QueAkAQSilcey/E/2rh/SSl3ReGZH5sBMxWra9LfdgkYc
qAdLBn1Nb+zRmSGCpILDm9/WMEKR3vaHiOOSDbrC4k7J7CeCtRX/eYTgR2PzlDB7RxtZwUOZTeqg
LPoh7fm0Q+8tDAzVlXKpZba7Kp4/fvgjXBxtBL7YwpXBcQJ9B7BPSbHfwHvyozro7sFqbdbDDfu4
lrHnXu80xH7H3j5ShQmFP4tRGMjmzyaBShATYM/lBL2X7MMJaGs3hDyanNxA7jExKqCPkeTR1hZn
VUueYBTmg0eBC9qhHFZ/WlXpcK341kCJn0h1eyjX+r/R/5EOEudQboASLuzYVZSodBrkcQJAJqyt
8xSPnR3feM658GK/zNwc4S11tmegfs7/0rnvtOKusxHs7VEW0WXnkQtcZF6jpTiuRVMSnvz48CYp
bXvskEOds+wwNMpC3ge1OsP93oTpN85VVafahHCpIL1cEQSWikO6Qk4g8yk4Nn1Rv54De2Nvu5mp
F7jq4wRvMADiyDibL41Ql1QnDFnslCBkAVUsnqY/RNDB2lDTgvjPfUNCVUfau3cYBphLFfMiIMrB
Nvuln0AJSKpX3mo1RPN+IqEjrBEIJrBxJFva+OFzkvM5vzxcEd/pw5oJGw7JzMDo5CSht1zQOXR2
BuFaIDyXAPPoLL76HKEAkU2y4z7pxgVY+xBcK1eM6SaqiPe0ENQPYHC+LXE7Ei8bkrL6soKOB5ng
OqkUbGjyQW3E/FBfsxcCWSidAcoFXgXNoPZuZ8q2baG/ENpBwpbUCN7JBIQhXy9NLGgp0tbbbNb9
syVGpc+BGvNXxCA0XrJcIIjcm6dD3l9fZsBE4sJJPscGC9tpR+gxL4V/BczdkYEfJm2HF8lvhIyz
cJfyAFwvcEKporFdUd7hlTN9XyIlXojCBNnKwG0XOMGwAx65rSs8BwykT76dnid1CcnikQ37+TvI
0MjNSxGBuj09kY6Fa7FIf7Tt9Dqo2iL4bK2RFn/7iXWDWx3OyFYvXCqdp6qKYKeEtfX1H/o3h8YP
HnMmJeSKV+55pQCXUP0yipT1gK3vsxpeGA1vVI/AM7BQfrA/Wb2CGtjXJ7qLCfejpEa6l5/WLA7b
aOGqE+6lg+r46pZSlNd9rXDvKrejvMf1gn7NBp98dVkaL/iM/X2qeVK+QqvTq9g+dX9x5QT1ZcHB
R8WZ4yhvJHKKgSEhpfFn0sS9gSj/q4vcArhs8Rfht+SPn/3r44QuxuUXW251wxoWmOLiOHgeV3fs
AShzQd2/qirDy4JGiOuWzRf6xhR5lVGddRpXfh0+Hz69MDOOf3qbV69YTbhXGWMzeegzQCstnM3p
LlGGnZRNhM3sYOidyYTO6EHds04Cv4AGntCyulYwc771FcQ1jipKAQGxFgdN+5m+6O99qqrpmQax
9cSYvzpXsokkhf41Q0T4LUGPYx8tux9pw8wtQCYWOTbwOE/Swin3KbODM0mWhXdMjMzDLoT++zSK
JCVwnD0X/8XOur/nQ2YFWyVTEVtfrMR8w581qwf6CjVolOCDoPIbBjH8cYdGrK8xy8QRxrC01BtV
p8vZTA525MdjeTKA/923xD9Pvxe7BLTRXFFXcXU/YrZp5Yd9tHkonGkQ+Rlgw13XJnQ7tI9SkXYj
b3ag13RIS5pDwLvUDr/VJw+teT8Bkb+bILzweGfR69DfJgw9bEy2HTpdgDV/q/dS7pMSn/LulZwv
yIRhvDlcbOy5vl3o95OWXOWVJTRpQuos6aGemYKKHq8LfGLP2krwXv+UVFURQSMndC5eBQ/Wokt5
E8MYBvPN6AcJ+M57wPNEoyZ5817s7d33CPW3dkfO41MrCFYnzDrZPT/vECoITyYYMnscplOh6eQT
xMu1GELVk+NVE/Jz3wLjEQ6tbbsaEoVvggyuuIkmnbTzhglP0QCicRsKWHkURqm4pRCuXDw6NDmk
J6yoBoibpRjLppkvmGpVjwqZRJL2VrnWIKcig6jFvP3xNgUNeCdiaSbBfY7UM6FOnnkhM1fyhSp7
Bf0RRxI85VaaG+bYXlq49zoGwRpF84b370IwPFheYOdh/Ob3/w77RjtViRqWAUuA9ie8rKiIaLAs
a5hjxUJquQQoWsTJF+A9nC8h1Gi4ACu9qwTaj4DOErIS79pppm2GiaJRBAVNrFc44FS8x+hZrbTc
HPVAkXwbCEezpGVN8zDQqg62Gt9nJwfwQHa3E3ZRqeNV4IDJa1L2J+M3iEWc7T+t3ncfoq/mtrHR
xCw93imYwXMl1FJt+OBKHvXtym7SepvcTr/fBhecz7wgOJNbrMZxR/vGu4hBfikpktAZYX77Iq5I
XoUB97b92eQpWWDSMmQlYE4dHadl7EaElNZNN9IXfSphM1AmxqGmuEij4IFPFGSI0z/07VPk+JSD
xlzvtUg7mBzx6b/tpENnOuP1ciKITXHfu/gyUQ4KmEZsXQntFpw8d/18WLm/UrtEUq9Q6z5UeqLQ
xDKnIbZ6giwEsXT1VsAhGtqRFBckC7kwTeGYPPHvpumT2YmxhsLhPGepJ5lvy4uHqCxbL6YDZwY+
UBgFAkdKw+HtbQ+QA3N3R8DE6sfTzweHRwRYKaBrnxAo4NH+/Da+A4rtIcPgkUQcqfIL9wWwA3OY
xCcgmN/wk2ZeB6jG5KOhV8b40KInfojMx8pAIenM1Ub6fLqvflKdjBbGyiY756KOmyQsuwnTzB9C
ZVxDCHHiUV3bCgr4DeKLjeN+OQvFOtGifXl/FUuK27gDkHNCmwBvdyF2tCFiLidASBBX8aaE8oQK
Kt1p5d8pYGiXUBO3K1BNySQDN4KnLk+3CfBk3EEylzCLj6S/4DQxou9ojR/YsVUjn47hA/YCFaJF
Y2vsbR5bdNr0lWAigFjuUrGDVi14gDWjMNP9rufLhtPW4Pdhdxe1IbIx6+qjYRozv9RldRus+xfP
55Wb3ap+0mJllmWw1iXsCr+wInslNG3D7RvCGeo+443aHy/Ef5ieT/vhc0mHQyQZ1nDDn3HuBGV3
PxNsrUp9jCXCds+eGR2yXSDkl4ZnrVPw4gwZM3jCQbwV3R2uf+wZEiLmX4wvOtR2ptF5O3mHgL2/
BnBpCFaM2pCxd99CZdJgBDFXR3bYXBJIwLmstBF7oMsKQ2YTxi3DJGOTE/bI2yE5kXw90VW++4Bq
vOPLSKOGuMldAKUdqqZZz5RcJ8MeqZ6MDZa/AaJ2C7Nq09y+TNJ1H8FmFtqX80pjqGnlUsOxvcqW
uJ5sDxftLO5Y4TC+RJdtUJHtg0Ore+VaJklSpuw0zmwFGiHUHIebN+ngQGiknPp0YZt8UBFA7/WH
hvqqnZFkB5sYqdIsOEgZnFU/L+C6Y4Wcy2GKRlVGsH1U5jBiyNNiQX0oRx4MaN1RNDKN4+2gJzv/
tWyfZP3pTg6SusngNG40ZGRcJWnKA0rEaa9kazyMRNwpot8PoHj/WndJL+noyuRjqSRZv3gVLgee
uPiiRXLfE6lsgm+kZ4ShZZLlZVmOB12R2uLkRe0C+a7rOSQjv6UJr6onjRaVBCqJsNTiN5K5BBoH
fHCfbTSmxFtPJjnlmW7JJ+wYGL+qLzmCgus1E3rcIGj0wH47qSHrLub5PBr6UNiYv3fi5AqOyCbc
pGE8hdIekLonyK8czRLXQOOin86J7uvPyOt2d9qcWASv0XKfAoTbvXY43rBu9UQfU7xiLRaOouo0
pRPT+NlaD8HIailNNGoqS8omG1LDxXZWCydIK9t77mx/YW9lukps/rvQwulpFNq35l/7Q/5lDbyQ
t7+dMKMWrzcU+Mg/k4Bwmnt5TeTQomdcIWLubuKnDbInJ5BWWDhajKT6QKVyHDX5KQ2jou5MjgLv
bHL0mYpVFJZYtINUKpomp/xvlAcUi34GOS0YnONRqZtVvQz/iBKuza/jaol3RLdQr3rN8AFcN+e7
fg2tNKBzONcpTako8EWKQ0gn0oFO66YFnChaQk489YfA2KmeD8zr+K93qEtsFKGtL4NdAqfAhbFZ
/5Oz8rdPA3YzLRRfB9rC8txy/zBllVi/4lGGcjGKQHZvdPDMqgey9R400Yzf+8YVme217LfDKAH8
4k9GX4NNXoXyJU+MewQpp2FLgEbQcUV6HvK9MsCs0QU3rb3+k8LcZj4fBbVuN81P9v7BDMApvhdD
Bb5kmlrPfYtu/hJcVx/hFXCxZknVx02qBpsbuVQ7x1EGDYW5zbwRu53azQYCbiIu3QSpRfLmwoS7
YsOeLgBwBvD8k03dEXxX1IITufNqQhNNk/UTk8kEyuDK6pF9iKs0KAw6fdvcB3NppRKQ3zJjQCWQ
vah1gVkPPW//2HRPXUOOWFPEuxHgNtJ0EuvFtZof7v/AyybGZbfVZ4jq7Mm7CeZNYgIb3w9KpIGP
3I1lILj3iVBuXcXjG2usd/4jc1bU4sF/b6WlFsDg3TWvdGdWdlc+kx4a+Eq9ZgDOwIORQjGHDJDe
AukOUf4pz7WYAUoN63QHO9GwPa/xjtLHzL9U0RGz4MQ1Bj4nmKKwIWnsLc+Qqdrm/fiWxPTdrcTj
UUu4YA3qI/XZUNWKTRkcx7/WRAS5pJg9+rX2PY/KyKPHsEKKp07/AAsMcFL/pgZQf+Hp/s74FPLF
0dvPPTtF5L0JYyU33Wk2LMfaQGCvCE+v4tv5rytyLFvIUvtzuoEpoSbcPu1DRCeUfcm8HdQAT9iw
+C01h62Q59lYoeJIWM8nLjleqo7EvoUq/7+QibiFcpB96XkKx0lSs5/Cuhfgd/7umStCl7K+lfXZ
Dm8cmcjQf7mHbOLnB9Wnj9v8HPWE6p//gE4cRhgq6noAf2nzB+fRkieq8cq4NS8qzgpUe/1idmlw
3blOwCyzAvFlMpsM2DMmpfcQCWN7p3UD19quczO/GioVom/5mXSgZwZdQ2AGE8O5Mz7pf27HC3go
B02k7xYFtfMIm1ePtOrVUeSDRpVafalaYJaN9NF0XqWS9PlfueN1jcHY3SUwDacCB/gDnx7czTAt
46k4hF6LVoum9bmL2FGVw7kJm3lh+enRX23eXB347ZSTQpLTPvgo0AW0Ad+3YcpKvveqiHWGxOjY
K7bxthhPrbtZKBUr8+M8gVOiiP4qeZctFXkdBi+p4FQRFUuFbKQnDr2n+835anuKa3UnxzsL6Iis
YPeE+D+P3uIuE+FtsNWj9LcvRyV+6SfwPjhMJCcQ+NHVxxyRziv3SHDZX826bSv8Ke5TkAefrmTf
1Z9tK0pAetY5ixm6QQG7irhMJ+uYoDit2LyqXOfFXQIb66KqQPIphIqBhHqxxT3ZJnATj2iRUlFQ
I2M618fe1S+ThoZX3g7ZoJPUZr5d6SSMhsp1DK1kgMR1rCbxOjkn6+K4vPGAO8VIzLqHO6oUvzZd
WLO6Vu/VoRdLIBiYw6V1Mq+tftPiuK9LfPxVAUOpMEaj1UX77YjiEVE4co725o4yWaH9poXFrpqk
vh7fjSxNyEO66HXX72XDi2uXdgiYdXMtjiC7KsB++z+1ZMpkzb8XSPqymfZw4kGeZGtuiSPrg0Tt
Sg/U/Ksf9ubpI94BIAnYh2Bk5tgJvTzhES5aXppj17PXPwTlTqGm7lYxEsXeseXQ3unM9ZuoWnbC
PmHHjdfys80jr+K8xhi/50zDuH8JUxCGr0Z1S3thiwKyrQ9kxf/Clrm+upPuobI2hOjsdeJS6wn+
r1eaGTsga4yE/S91gPWeP/cJJk/W3KRE5NPos02OcVbFfcxWeY2KaihI1onFIhfv8ViYV7g9ZE0D
ZqJbF5OtbnFdC6GorhpF7rgTml4Ridj51pAXVSoJ9pl5wR6PjOu/8l0jPx8OoPH9hlBmOql1zWfQ
0G7gyQvlpag9Daw/ANa13BTcJAuKGgLlQK5lhRxOI5qz2fNBHbBRx7GzIjxthgjX3ls3gzFhvwcd
SgwTQ2N2z0uYRul2pVZ5DrxWKU438sZRl1DM6M9uJZ9YzeorWY0V8ylFHtbuD8rf0xgmYBeOMw8c
km5inPzffQOyEwrf2KErldSbGQei9w3fJg+veFjF4l8BSHodq41ybOP0imUiRZ6Fvs2JoQwIB8yj
/dsPLqZBfqXKH90tyQ1HmqUQeWFDs2NM3FE5vfWrnMBUgSSUq62Ir+YB7JHEnqi6Kksobn4WjbQN
zdHMOROEFMx6hVUdC9nap5sua/j1u1zGYi3K6W6saLLf38ZFh4142zIYw6PUS0FNB6lU60aBOKz7
+lBFvJrvjon018zD/+ri0c9jqyPz8qFnYKbjM0reiCFTOdejHAimNmrvamvlKiZNJH6A1i+B6a8m
s5hZ0184dnhcLWtcDbpOY+zIIZcyxnkcCqoQdVoSI4+uo5nAsy5liXbl1Anz3X9YZk+5lGYkY/cL
cUWiTHIyRqAEkxsKbtj3k+m7R222piGrUYO6kSwxrXnEWGTKrn3YX9VZiZlv5bDJhrGTWQ4lhZSY
rQXxP3DYugPJhWCvwJA+oy1z09mMtda/clx2L+T88bPY6O9tYCOzo2JTPGdEA37E2fLs9rjy9afD
hgPqHjoKgOU7IvQJnn9UtElHas7XlNkxaX8hWIavAOA9Z9uhRtoKUXfIE3NNtUK+yE4JIPgAi5Wi
1tZoI+iUuwWCrMd1n3cjdDtx9wv+HJADWa52oHr/rvsWqtg5SpWKQ2HNX15YdpRFzpQrRZItMcuw
OOBlJmRTuwgz7DFU9/kG9+iSKDtpFU5CPXb8/lXQLDLvwdIsszmvLmMxdCSMesyFQqF14IRHgKJl
au7Ckb7xDAmiiG53a/dAWAOjKEH8gHSDQsUvqtoj4Kl737fgC1StLhkUXxAhukTzJ32sceKgeRA3
gxCcBpCup4bCAVflIaNCKpa0Dz8di+TCpuGxv/7EairdCd4lwVdrywg1QbcIZhzf1jpShghqol5i
sCXI3f0us94RMuVI3xuFZmiHiNDjAYzcNogaa9hXG0dBL742E8sOLj5d6N/A+CdeKw7ATa/6M+Ww
l8TORnQ/tes1iHdMRxTPYXE1BeYalySoVqMlJVClKdkeXTEE9ZzhCSrt3dDx9Hl3hAVUe8SiC6g1
ECxNmaTDvi2DfmnOcUXlsoIC95ilSkjfIa0vEvFR4unkxxXiUZHexJVhAfwvp6kFPUgdqLrnGgLo
19bdk2AuLVJo01JDyVHOB2F1CNXU3tth10vV0kWDMmBd/W6KPzfnIuRxQTxwpfnJmuR4OvWZANXY
EKyIwlBItSJr+HrfboabR8IUM3yyDDypu67sMTPvzFyloOqC98GF9KjcyCq+jrB65x5YbJPjUCC4
asFrl/8+E07FYLD5o1EA018hCxaolmr8vGie+LSCANXVFKkRuFop3Wh1lVi7CnCn8AkJV2NSM9mK
9h4rUkm5AlkEtdc5x6XgkTNLHgBRZww50EdAoZQuKqj7gjBaqOQANZAx8lPKdeRFQeEeEF/EfHdK
1lNxLq9vDN3cXpdhdFJUlVV2T7kcBIPezfjRbxGU0FCXVVBgbYat23DDij0If7A4iAVWl/L6fsMy
hxL5BHwUscJpsxZRHSbZaJUYnr0NbLHxbcxttfzDoNa7tn4Bwf4F1vn+u5/mvHMUEc+tjfwuDDzm
X9tRWlBw5U83Jw11uwC7bd6i/N4fkMU5u1zCszrb1W8rbwZw/+JdfquUcaWZxLvdKIOime2NsN1n
7Edmf63iQimbC13MRydAyEw0kBhx+UsnN707FuN2XF+ervmxxP2FqFEMCp348OhCGRwS1K/XLw88
KVqK/SiD9pJY9met1dLt+MoHqJj5/9qpROlbVRte8D+KMwscI5aC4fyHN11/qMb8WgXermE3D6Gc
jD4dg2PLMxo6gbz5Q0PUJ09pBzZvAtu6dWi/4QepgRdBuzmc3D/XivQ5F+GC9OiaUHyLRLxBO3pY
hSYSaJKqNtss/qvrduXVSmnC8P/Q8m0KN8jV0dddGwy/DzYqwU02KJUEhdPdnmWs3QX6z6RKdKeu
IVQRAT9BStDZYhnoWjMmxd7GWEtlt/3sT2JBsr3qS+AcolgZODNdilhRZnM0AMmzDG5dDXeI66S/
V28O7ir70G29G83NVQ1uAI0SkZs3Mw/OEgF5EidP3D3TOqyaZRNm7tuV8mQ95BMXayPJ0ht9ALSZ
1bnfSOJChf4YLIu74Q9ZpDbt3WPevKpr/OZpuoOl12ExLhfpXkOrMO56oy5QDZIkyTc/YFhf9q+y
fci92CHh1nlFfT9T39LuOouEw3B5H6Clb0AF5aSDKJ+ktY+/AKaK/KhI0cLVpI+29Frw1MYrTEXE
LIwrbLDyTTlnIuHrmyvtYLQrhRiU23RlyeIreuvi+AqsGvx4YiC4P1Pg8DOgXplMUmFT6u2h1eDj
4mEGKgggz3h4ZAPPK3oEKn8AtEdv1VQTMThluTgLNJLlpXSSY7UQtebE3xj79gCCBBH+VDoY+JHb
S/9koGR+0jTYQAi3+CTGUcri2+fZaSwj+pHhfqJ062InWy5GeGZ+fxrGM34XAkOcBdFZIG4qtPZw
naI/k3QTVk0ETme7JOyovYteR0uSbuDU8hi/UGgrKBF9DDHG0tm9VEn+gqTDR5tn7jW1UjIlH/ch
GgEellb9DWIBvN2xaao4NKnasIba0VkJSnATCGOrlJHXTvj3Lj5grpqvwtQNwd/0P9SHrhDnqlus
C2OgfVjoV2jnsxarRvMQyRzs9EvyBgLMjrTM3kXFiSOO0nTsRBtwBhzpAzHVCK/ZEHc4IRXKtTEj
jRTaaiVVUDXgGuivZKGOONxhKQjEV1zhCy7Ti1xNTUZUEFscZhRIzyr0v5Ukibb7R183eWCxmrW4
jMJEj/i7Qar0qZZudN6dv1Zh18Fiy10JkIXRJzDyIsUGrZy5u1FZ9GHKc6Il1EdJ+RtNA0ml5AZW
pv6H5F5OCMDOnUeIy3EQdF5RU8fQsUhRSjo28lLZhrw6V1tBd7W7GgfasI7Lr3FUZQUDSq7DGXkd
on02Ffk3VpTceTFSDmxVjEJMxhaMZLqJa9wkqRsCqMxZQHa/lpxPL/Fj39/Kw/96bw4u3RAm/C8F
9cy0gN0TxsIsgFdQzzBdjWBwHLsn5y/0P3WTy4ZwrW55eMq8dmj3Ym8DSDAKuivVYM+BcpE9r0sP
7dxHLqKbrbXjlBNjkn72sFVl2OrjbfBXzWrBd3SCEBmxG1YF3TIjhDFW7F9A7LQFpMDdWzFtMGTe
TpGAbYdD1xbLNtpTJjCkLM+09H9J4NLw5iFYMcM49ugsECYyAe8Z7KAk6VYxKVX2ltZ9I4CuRSTU
M4jiAs2DgPbrBL0lceiS46BE4BkmeWbxvFa95NPdEbbL9RXEkkUzJeTk5Ma8aBoBhU7v9RhRDYZz
Wq/BsSmkqo+I4bs5MewanmwhdzDQ6ERhJ1pfPcmrkR+ThF5CChXmX9cX+jY+eUhhRRHYW6eXm5SS
CcR6qgzyqroP32+3mc7P3oBNTqO5AQpic8rol/9cyUojPcizqABcDfW6zr3sDM5mbh/jJOol+4JL
ZUqOKDiemk7Xzk8llWmW8nDMVfCYPoOOU6xnXR3iRTyt0y39ysqp7AhJQdoDy5HxEjNRvifcfvmk
4uW5N6dElwBF7b7mqPZKtRPhh5JoBFMFXvaGOmFIComjXNdGROC1LmtuIgWnbYkuP96FTGgTB1w9
+UeUj9VrV+f7sDvoR5KZiytT8HuWZsPFbTLFZKaI92f+FngV1DA8frTaQl0x9mbu11fa+i4eAvio
d4Ekl3MYTGVQBNvqLoFI/ho9gxwybeiOFmqvqJcMze93F0P9G1UA4tlMzPZSgASakZSKerC/3H4o
+D+HyvvrzWqU9XJaYDlAfiEW4pTjHXF4Xrc61vE5TGXYx+F0jDg09C6cTD8XSPDkJmOT/8+zIzH4
yjku+ayYjczCWw5gTVZhTT5G5UqRURlkXsHlycdjry+ZhWO5K1kphGZX81r74eNut8TQUhi7CDVR
tTuVhepPIE5qoDba0B2tgUINu8QbtyRkUSdtF1SJJSprFu+kYejRo0PAfKE1eMDl1CpZ1QmNl546
JJZ7S7FUwAdFYVU2l3BcFdnL920kG4u4RSEvVo2Lbv41aFP9Aru7LGtj0pSsyDd9x9zjUnOQkC29
VhSYIwZRpYpjvd+fPaESKUrM269gWCCd/YZH/wzeIMRYAY2akGw9XzhJs/wIaEQA8aOw8/8LhJQj
K0RqS44cdaI0Q+JkyC2GSuF0by5Y5rvVvxfW2YrrCl+5iWMWR7hSKCy75rwlGtjFFJIJ1pChioeQ
4slJu/tYgRLNL0Yj9KWl5BQ2Msbo2uMV6TibNAymhH+GPxjOsSePv9rgNKgISG/P7+WoU+kdDHet
hC5QKHcSR3cJIKLObTcUmFob3m0Djvi0zpnsHbyAtVevNGkKqrh4lc7+g6qNzH86mUjI2LqbW/X5
34VnOiHpG3Olr6Ff2lyX9iO2oqsbY4UV0k3UkJFZCEMeou1uu+4E1LTVWVkk0f0mLOX0oXI51Sc5
228IzRtnHb/ybWa3wPeQDkU8qQHshhsDGDaSVYMODLiylqhYBHMzwwoZe9SommpLcBLuNKPtrvMq
/IVPoniqIIFCFGzq3iWidvdvsc6nlBedzCXxqg6Wzwzc95V9kk7ti33a7kkPOSZ4pagewjV7Wpeq
y7pnwUhSP6uum025CXwE/CDkr/9FU7KGBkluq/5HTF6rFM6QSQ0T3N4G7+yXLee9x0XrEhsNP8as
iiUSlWMb9OHrCrAEDJNKc2gU9Mt9iNy1hIt5U36PaG5NIcxyWX6noJ6fdetulh3Vc0YYW/HKpLjt
vyyArR3HBdHpfrQauiQ1QozS/T1TClefK7kH2Jn+sxn7A252H+lRKimtrijr5z6o4r8QXhLck+5+
s/zqJttP0F8/gAli6Ue3lOIfbotqfdKOemc8C8zaRc12VGamABp3pVxZK4l+49XwhSJ42bzn4RR8
koVN76xAE0klO1B3AhyEI98VreketyNJrC27Jzb2mVy5CYw/k1KdxbiDdwWyRuOk9gZ70TKhFS3L
HL7WQesf1K04yz/5wHCY5gLQHX5a9zxYjUTJ7LJWE7sqFHq8usNfnasiwh0Ki5yy9bDRQn81bgjH
7qTs/7djAib0bwHJOtv8B4yeJl7ajyijxA2mnYm8BvY0ZVF9GPG80BK07f7LfGx70IybW8vhfFtg
3D1NSjLTUNj92gnNp0t40r2ati5q0B6ezVlAZzaS5mtDwlaQMME2aoojMlow39pzxtKnorhO4M+r
vJ+FW4Dpl/DDdI8Aq54kB+Tlp2n9SRetv8FQS4ptthh3vJjHBp5foBZigyH1vmRdjkEPqU64tsNQ
2zc9invoNgY2YgbSXEjESzZyE/tvu/qPP31Ng8hMFVnumcuppE944lXDVZ5HXXluyTdmJhJCF/yo
e544RLtVqE1HrIhdW4nWfqQPZd1px1WYo1UT16+cs9pvis64tYpG+8K+TKu+OMHyDA7nEw4JMMQd
1f1CTNGyx0DmqXnTfH2737MZdFudyP6UnEt6kihVJ3cTyP4yqGov51qn1GZWxsd2jdsRyhqS28CQ
oTY7rI+KjALBSiFU63m85YzQtqHQns/Melw2wihsMLLS7WFXGmoKj8m62JXaC5E/ZMsZBTnhkbnX
uFaIJ7B+OsAutGH+HrOB+D8/sRjrYkjMIUYBhVDYj/5QebUVwp3O/FmDglT2ZsFTEcTqNDUITDmq
bgz4BtLSaxG5OFAvcW/lgWJ2miGMo5JOFVpKmLzqBHKyq96OTtMq95xqCoGdC2qORgjVvV9RH1DP
Kf8n257doCqKCzjBGD0Rhb6ppXdIBQxr5VdcrX0iJ7WBQyQvaLCQf7tlqRRAQyPlxh8PosUKEcDH
A23cEVcNuj1PF7hPMDGuzbnbeWygn5DdTzxq9Epof1+gJuOvegeyaUe8kdMdzEbQih8iZt/dAR7Y
649ZMb0KfhIlo4qOdbg38K2zKPnO7uf3ncDD93pdydQtesU4Fu1QXuZ48V3Bj5o5WDEAEkVzgeKA
iwx9LSFf6uVGk0UgYNYsWgdtCHDiDwy9U/GTh3W69F/xYMrOhi8K80wfb5p2DGaehlxIjk5dueiH
DBjBtkFlwXWOEVVN+FC6dj7X7Sk2MlHiBKqo3gn6TY+KHkU8hRiUtK1EHSMKf0+iXwyoogu/y7UW
+FW7PbZldrFqVp8K2r7XanCLSN/Kp4SY2RPoB96HWkOFBas/x1raFx+6NNtMYmt3VeKCnhNulUqV
tsDnsn6yrxXJ3EdJopiRJjJCBvJSrBmSU2bAtrSR3MFtz1ivzAFnpAxWqcoOqS9fmCqGJEX9Nu1m
ZuQ+NKJIcLy/0kHkkmMvk46LPMbiN2yfplg2LaVOr7LDowNJ+Hy8l/PQlLMPA1SLttH5Y2bZPJcH
lgrQGNXgAla2nOtD3wS5WFxiocV12yaMkikaqYUGPPt8PRzt17yNXjXE+5Kh0hKN57nVKKOZ4Uri
fEUIRFu4uaF4oNhzJ/LoBxZitTj3IvUt2NFIt/pv/HMeK7e4GTUdDan0ri0N4voZfcr03eW+G4Q9
aW5ymwcow7jN125XpsPIetzsHT3BCpR7v/I7YV9D5t3kLEbXgvYt2Wso05sShveYJDb0TYjTd68b
2cDfiVgGgnJU10QuotJ8YAGzHEfUb4LQboDOE78FIwtL04dticREMZViSlSBQHwCUCELxnebVjJj
2vvkUePJlQHoo5RN/ms6zW1GqI71FdBMdiYnKn+lZZTE+eCI9fy9Cfk2jiipkDdhSAvovNjnhQ1D
XVGBvFl5L1S9HLdxyP6L5BH60bb9zQsv1yS0+L9yBASlPFIj33bCA5f0vs7rb2klIPAmdsBgvD7z
oDiDAGQFTHpopaKmRQB+RkRraE1kdF7VBByikdf2DSi1Dpz0o2ng66EP6A+Ei1QhxGxPwMtbUtDz
BQUe/k3nnF1eKcyFU2EnSUectjy1uafjPNzCDm1Mf6YJoE5UWmaDl2AuKS/bXXwFaMcVcUfSgXYY
xRiEfFMrlpLRCyRORV10+1QaqWRz1w/7gvUa152cWsBbgQC4sFe02LKGJ4okID8/56O0a5T/oHsu
TkpKc7TJVjw61xgOQ+chyB+wWPhIzMASKeKWh662aDygXFM1ehqs6gNqvgYDMP5tj2OrQCxjNsaW
1bWpSP6ixfVgqv/cuWftAVsCv+tw3YihPUsXOrznkCr+pN7leIw8RekV39BHZCiHZRQHwptPXppy
tBc785xHyKvT60jvo2uCeZib20psM4HV+wDIswiRvNG+pDFbcfdDsDQYO5S9bZhMFFK2bfIdIiUA
mn1N/By6tr+XngAUiiKf3bbvh5cYnCpMVCrNkvaD6+3E/DIHU+Is5TvLA05ES6bo2QMzhXLrGq8S
cghb+IsE7vKeRih9P+sFsgMvE5FazgglYl4+WkWBxiH4mkwChiGHZE7jvWavZCtAghUz5h9nleQH
p6yjUqckP+Quro/cDyRHn+pKTXujtyy1dX07SbqRksFH5AL+QZjzTd1/81xPtdITCqrAOlTeaQCm
l3/QlanodEN4kNXByXMhZ5ALbZ/zyjBB3ZoRTziPS9NtMkGDUp5nRogZAfK3CZGHorK817M4lxdo
qjOOBfQMIMQZwRdVueM7Nh8ctjRxQ2/HHJtHLkaVxLxHu9jJDGYw7exHxWMViuKeQ6vb/MWlqTJu
1y7Q20MPga2UbFLSizCVSQwlfUK17hrjf6KiGD1lU+6cm7HfAGdFecTbV7lZdJP0C/Cxsyo8IV9e
bRqNpCajXwFgs8FpAjI3PF1DiSy2ktOqsjw2cRhEeMXDhjB8OBxtwienw24+GNgGDM+4ICC+6O11
HxHBsx5xddvQu90HnTHmy8dhtGG1Iwo0UXSn9IzImGr3znu2NgtnT9h/Op9IhXrhbQLNKN6J0RQb
U9OlzBzGUACO8fq+TzrVqQk5DyGiNE/x887cJKvpDc8TSNHmv4i2s082i5Gd6GT1ajzY/UtVa9PW
E7yR47bYCMRqBTTIs1pvrC93LiuDmnXPzYuCrJmug3fQgrBXSKODfdTLgOHfUlAXNsGz1Lk7QiBw
HErrpF0eQj9i42AOUlz6c61mNhrmInw1asWrdf2fhMcg6x/2ark5xLWbFkiO23Jc8wtuAA+5+H9U
S1jLmauCnT8YuFt6lpZknSj4hjA+FwH+gdRBrdof2xRxdww0glgyc5uhIdcyCn7kJXdtZh66PxaD
1YbFpkLxBpKY0+W7k8RdsrlDQNaFc8i5xhPuAwwynGhntLiSDDh+X+D7IRd0DsFB20UM8oSqXQQA
y+uqdsKgVLitf5IODHjuttEfcsmHfp8BMIVFN47Ph8yyw2UzleGfHrZ4goRCRU4LieDWrjgHkxkY
9XowPuiHsiS6PS1GRjojR7ShPnOftU+2+PPYTLAQDzmRoTi6Yf/iWjlxl/07e23TRfIv93FfpRYo
yVxOLUE7rE2HUCsaHwGkC+7Drq3YWKmMkQJTTdRCems3IHeE3hElt+SVq9eLWHhjlBY+C5Jja3Et
nRaE7bL+dBS88UNeLTtHww93TmLYi0X6W7VE7BZ8CUAi6szkLzo2pC45qJZc3Hm44B9ciR5mxZmH
EfEwZHuHt+44Vhj/Kc5YwSShKW6P8Cz+q+QYlo7zdmxnGcs5zJtcyXOj11EJHnpWoHNFAuBmQs18
JsY3hEq1ZFbCXxi+xeI/FGauwbgqmmeNiXs8FNkkxFhy/zboNe2HLfqfj3BwspIWJw7ZVSu3gq3F
WiIYMNk/GqhZti3W3jUiITU0Kky/DawwxeABcLoUQ7u13Ao8f8CQv+WS2By4qC0stMCcpLEP3shW
0MeKuxDP4zpvm0Vl8DpJ7cBdhlcj04pBHU5WyP8qLVDMpAUu10VuyRs8g02qjUvFxIDkGBAR38hs
plt2DZ6u8F9x3Ttzh4AUhzB+M4dM/36gCDUdcKmtSFXJdf/kaEtKV8qz/qhUMxtSOZm19DCjDg2z
cxI33zUzr0+04761kky1chpzk8r3W4Il2lopOlZEnXthUYDMckVcQgJU69sM+li4EmvmJbKd9V5A
6+LPB21XPp7m3B8S1hfYL0nuOS2GCUecnJCRBct/R45dlBolA/W4e6yIbH6poUdYLTRxjlbQEy8E
Hxpobd4brWTf2buCQC0iQTk3+AOHBBqczlFtt5TNVNLEEQChQ0T9JLe93e1jveMQRosc3PffpZhF
mJbVxuZGn+absGiP+UeHQJdEOnC4aghvr+hKfG55NqB1OjbG9BcH3PPL+aBP1mMLsTEwqVm3fgme
gPw4XfM/p25mvX11FQLUMzg4TPNQXZgs+HT7Q7jEX+6bfIY2JvYEHJwTldpSU9iUec+nLQpAfa5n
7u+au0sSL41vwplchVFJ/jvWOL9HHbUVozF4H5muqF9TuycVldJqeWZhNT84OA+1kzpW2iNqAdtb
OkVpBd1eWK1aWkBKgNKQFht67NJU3yQH1maYnu2U60sWf/JKQrrjcIais80wOu4TLsR5ypNo9F+7
OOuyo6FwFIuGBpFShoNkGxa9k0Y7m9VfRwf0MV9A3gSPDH2mwlAyjni/FQd0JenHrZPRDMzgEDcK
2y/5BJfzOPKfz6zLRq/XL0xeGFf8/OLrJUUnQ61ZSgwHZUoXRPO3NPCCQOjwLveVmMO7uW7Hz0LP
RAH1N48kRiGJa158nuwsTrP056keUv+VemV2jlP+uJ4ecvq2SL5HZRGi+GKfXOFSzQxMKHhj3vWW
mfTb97cIgGse7zgIJnYg38ztkhVXgTJCLWTtT7DOE29NWCbi8uREfKi/UI9ySeG1TvIwLR9HKxH6
egoOl7wfNAuge1p4fnTYMfHvGAaola6orGbzWE4Pe3wRkIAscAUfWqif5hJ3oeq9WH1C5YcuLVL1
FyT3bvwIklzT1SD42MR/iqOWhyFAeM/J9Rd3jQBfDOtYI0tf5ihiUVxgm2tDDBZ671NgWOxGqhrI
1RIKD2dR0nObOmQNPhqlB1rM2bpBUPsKhdkXT3lh6MGnfRdj6S9ZNnbvbFj764obYmBHgYjGRBFz
rhEIRxbTzvdc40nvRvgg2MBP0zlhP9S5zhXmcweqSKzG6lEnbKqQsw5rLbGFNtqss5l97tkdt/jm
id2+6CNGGSNyz39Tg1fWvpZy+r8MhjXciFsFlt5TgGPCL+YzKbHL7MhGMRCP4eoKqoMZngFoZtcv
bJzQgZUlN/P5kcxbnHyEtRnnXPtQOobsV+SAgxCH9hJHKk8fIcl0QeCali2oMoZF9Tevb7AcWVlW
dgku/86MdEmU2eZDWcTjxXzPht7DZ3E5qpoz5cJsc1vmJeYbInI1gQmn5dBB33QYFJmioAfmXrLe
nSyU/jcc5jfMdIGALBGrtlsKG8EMAdieUN37dRGRd41UZSGM8TQzYvhSZuSLKPHpstot0fsW4XXz
j1vzqprm2k09AMuwPIgHTv2UO2W/IlyXq7z/gTFhE7ZjKCPzUHG5qK3IzXyVe+NhCGMel2XtyCFP
ZVqCu4jpWaRaKK8hvhclNRkVixV12G0jBJRGSkfzq78xUmtk6qsX29pWT88yFNhlLjnR8jTdm49W
ZrTmu+jmiUiKwofvfjJBFtelp0CwXvnIe9HLIcrr6IhISF8+mDRg5Ihu8y1Z28S5ATufweo8qp3s
Notam/ECU7KLVPE2hGDdzRgI5N21+wUdRPvamJMwhQ/aeEbJVZxw/xPbc3yHHC5xXImeMv5vMziA
j5aPcVQZUzotbiI45R27uh6JoHbeQgeOcTCv1QG3QK+MGNg3vJ4qhhMK1MwIB+HcIaY54Jn1+vXn
1ckYhmaojs5Nkzz5GIw6+Z3Mq6VFJw9STZHokvAu0iWHzqDaC2fxp/BHt6sxzRXy2kUfjDrtxmbV
Lvqg8ZWUecM+2UEc+UwpB/EFRWojzBZyC6BkEnU78KZqzyqFBPcm+HOraMA1dUmoM1YDdlp4ZcEJ
j61fZVDNou/1u7oXU/pjl9oDPplbEWGf46xKU+n54h1PtdDIXRxSLFvDX9LN14K17JjXhdQ0q5Aa
TjeF2/h18EdDuSl0MkR/l0l8nNedKIPMgnluaH9ZjbqI61TgxsnSEzr3Ti6kRRKxjqJHMIblYX57
iUoHBilbmkEgvtbu2fqrbiI1l3tyF/fJ+7t3tz9EXV+HaI1i/+KGPpbe5jjDkM4FMcloHSPDwNY0
3ZQJOyVPeEjtNR8QgyN4g92KF1sNf2ZrrUoeNH50dOgnZUxzDwg9MCDD3bXiqdZ97rnnUdxES+a2
3EqtyodlaNUvdXhYVJQ1B1YHon/vN71Hs+COuwdZAavySuBKTbbl/K5b3DxU4Sw4ed7PcQN4CWk/
fbVKHczT0C0BPK3mNtLc+s6txB0vOSe5NDnOLVwHkss1SMObyb8X7P1QZIlIfOdoqimGZOAby/lz
5jF/+VIDToCpovLrmfhOSeYuRT/lhaTqnK2mKCHaeUDdRD3v1PccS3rUcceyXkCIEsGMoV414sDf
sOuOgUEn/bhlH99X/oUF/QBGYCJgYeNvBsFbgmjC8XJBFSu5KG3dQoLjkPsDqACH6aK9O3vS3IqS
qeaq9v0m3xHl69WRisTJ7Q4cA4lqtPJc7yEX667lrZLj90NzReTAwEeb6dZYusrWV0qcYzosHK4d
NHeDY5LXaqdXQDuYTuFZTApWf8W9I/JSoFMdJmSnPB/dL5glpXMX82I0PAVk+X148Po6MI3ZVP7F
Fwiv764ehFt8bCkJEvBuY8DLF1aVyfkhgwzxZyBLtGsFM8vTBcRoXmtAEGRn7IxZ+gwDGBqPIRWR
kRuFLsZkau/j/kY9nB7HKBhaiFD5f0f4q6lw9QH68Us8BA2aVpSP/dLbSwliMDVFkSPvWXtCwT73
RRrjYxQmoN+gnSNUDtq3QYF9YJWE1x1magQWlzQ+SjanWfVjJ3mPpAOJe/QBvlh9y4RjaIBYwvGO
Fg3qDYUCrhIETN3NfUE42kNDIHYjUhoHd16tjcvtEJWOZ0hYbj8zz+0b/ZDWFxcWa/9YPJI0q/Ap
r2At9BdR3hdm82Hzj+KtxRvhx7wxF7XU8MBPsqG7i1PE2SDgrmEbL4+aTP2IjWzrmkvC++em2R5c
ngosmsnJNi4EhqPiy+jxyLxnqmVnFNZ/yK2hZ71Zj/jQ6K8uHPvE9uJgjmm7KFhsIAqN+VjbVsoU
sidFVYsQDU3xN0muYfVYp1S5C3eJLraFsD8G7u8Z8oI35ObthY4OaZCF/Yvz953tmFdrFFQHX9Fx
RRVElWYpxakkviP0f+YFYHg+E0cA6mABzLnZ1sAYycqAxQIifG8GSuB6XGyzNtSgdZAjNN5soiT2
LfcL/Ye1awrnX3MrOUnDlQCSLsYoyNccgCot3mSuuUHruGFFNN8iA7GOD/nYKOPMPaXfrzfCShOI
lRFb2CAzDlJcPQxFuQVUPteo+oDZKVVP1tNixs8HzXClDUguM8whAZXRitffzVWzg6PntYrvuxay
9LAX9qPaIy5ZquvckyOcKXKnw8VxsXXlTxWYctQMRsAuWdhN0669jtM5OQUccGTIH0cWOknflBxF
O3avTz+gQmibqI56OzO/CFULT9WxHNNV9Ij1HbihH+Rmt38IzDL04A3L/aJFTSwaiwakcdywbr3k
Nu3iSi2gxgMoz54Jmiacv3pM60ueM9aSr1JFhk+1SuQWM9SmBjP/rMOIDFjwdufUZSFZVGZuabGQ
BDRw65k9eF64lG8mmbroatkHOJjf5A4qY8AXLzAzR3blK23AY0ycuPca04SVFYKjPkpPskprlnkF
ek/dsp7MD+pVIN64d75mrhGwj2AWwSn9R0c/F9a1QhfLrRepf4lbZEWmbP69TuIWSpkjcZp/LmEK
EP65i9p1luzUPi/TS6QKVMNrLfeAXjY+/2dVRwDGyLPg0eXofIt2Mhkx2S7911sW0NiyeSIZTFWe
GuTXDYrye3RpKKSyDRvrPaySxUePeElclTPf2zfYL2UYPIlfOvHYVlTyHi7sWJ/k9BrYXZl0OwpC
+HL/FXivHa6/5SyHebUKmIh1QZStTuZ6lBdJyJIiP4RYLlsdPI7S5DjFhO0aeE1XAwD3lLcDR3YD
1Uf64LvlLDmNpnREieqIUmbioWNNWmmYEkOKnpkP5SjwozO3bl/0QbzoFssTiqXoY5IHzKE7oXUF
jRxJooHfCG8lKmPPCGBoL8VcEbhzF0eWgetqVo8meABSLq/C3LGtjXJgzCEyMJEiYp2YnTTjo685
A68dDSZ7kgJeTpV3RWRo+V292YQcVVwRuI4XF9RX0agvbzZKvNBJ5JH4v3mHFEtDnUGbSOsuisxP
BmhBQW1PVWx0hQYGK/sVapSeQs8TLSfIlckzjOeLVtOx6yqxOVgX2nLyR2/1S7+UhmQoqnLf3dWf
96H6j4Uf5oYP5dhO5PzAPGKmSnygoh/yQ8xPRc/xIk0q6AI5F3CRxCMgSX7hUrdTmUz9qxdJryRz
V2V/M5Q/WUjRDVFbJ+DqaV29LaMXVm6ifkbIzqTqds+iSHZ18J2z1KofYWmy15Xhu6U5mpgoEsyn
jhps2Uyg8HgFDA54jRtNKPCdkeMWwqOT8fBYQvufhRtmslMtV7qmMN4Af49D9dRObsPEl1U3vx8M
OntCtRLCHOsDv0/kU1FvSERjiH7WYq6zNkFucPqJ5TpqsQ/2GV4QbUAqzMgnj6KeDamEGXuUCQcK
p/qyQ209rDzNOY/Wut1y9ckuMPilJ9S72H7T/FHlTlKj6DQxeCx2D9BMXtvjffcWI72ly6MvWa9C
rwQOudRAgRhWJ1kiOxSFPvSx+3WTBX9alBWHgw3AQ/+qhVLZ+G/PTNFVSBTHhLTSGXmzhF+eLPSl
EQgiFsp0+ii/NUEHyyDD4jMJvLdEjGZG7NhhJLs2qLIzazLm8fOe4BctHYrPs58rc5BEyw66bjnR
0QLkSPV4UYH+wQCvqi0nDp+R45IXM58RVA0CPwBrjNAEbQapNq3Xdm7CYRQLpb5F38BBmnTGB+Uk
jPparddXAvgsYQwHKjPpOyW/HRupzT+THrTB3o+MdTHzIkQ43UXDswSmdr+DPoAVVRG3pSbUUer9
3FpsjvntHSHFbaLcyT+0vaiccXQijMvdvz008UUieOqaQqFCOb7dmSlMkv2y/MP8+vXd0PH6F97V
FrB4l2Cqqx1fgPIxWhzDCuwLWp4n+tO+yQJGltDxSONv8IQJKs9KvKh4q8oSvxoEdDAiFT/J5zYz
oba0PPGjz5TsF8eEcZjnY8CybCJ7t4FBy86hFi2ICQYSiCPrt/+cAX7OtT6GfkElt0+yBT4xC4L8
kEJkRrCppEBwJPG4xgLnZoe3g7QQ0YJULKLOQ1H0bylsnSZ+/gt0XAsjx5x2kUAa81hbSoqlXMdt
6eg3uEARtfKGtjajsvi4DVUT45YLDTcVqqH7a8vjedhhkdfXqCJU7QQm9d7J2uiUC0yPVOxr4miC
2tgyg1FCDh0/rbZFNX2WwBZoM7X6Zn4e39LO/fj1mQ48xUAOMEGLL01kpLd5TUqLp3lKLSomM/kO
ZAg2pW+ykNPJ8B/OlsmA0PvlQnc8566mYrG3bts9axELYPofPy7B7zljFYFsC4Ww4pEUAZ84BWcR
Infpku2dGjWpjTUwQvA4AoERlq0vuNuMyJvkTdyUpCzikL9108YPSbTmkK2Kogth/SyN1jJ+K/8J
Ezk3kjyKMs9gbLk/h9YvAh8XUbvO+KZgjlw2qLMrbRHqtsPE7Qu1+kCC+hzQVJ76eK7S4hkqdJ2g
8umhD/O4xOA0lAV3l1Gfps3550ZfEKHpupQXoA05VdUtDSFM4xtR1e2UZ+zANk1QncnOC1vJLfq9
kTHYkjR1+3peCUOqdcTCMM1SjusW+V7I2IwU2q3Ev7irVpxhgwag24Pxpko3YYgQKEUGTKBK4Lgl
LUpr/+jopiNYMw9wkripOwlO3LKoHvVdvqbfJlvxlKigxi0VbaOTBS6DgRZItlFIJ0XSHG2kB6GS
bJ7yBK0eAejWUsayqrMt82ZzpV4wnx0udrtT67FPHKKkT8BtHvrUk3JxzjApBQtCgaCAhqGzdjFT
BRH7LlswOjgOczXu+73L0Sa1JrDvlVAWBue8P5Vze9OsAkuuQvRQRWDuykDrHhsZUNN29883ws2L
6dXXYLJUdlntqMAt6LNdxa/IG5NC6AYdPebrqyNdPxuGANhQGtu9dGuy+Wzg3MceaJ+/UKvFJzr7
kVeLFk6wZO8J7w51HtxWdBbWzLjrtswzOYYuz3OtPLU0JhL2pzqiUQCgXngCWIfJC+b9Wpb+gQGo
NF31lFBvEycCrqKChlV7DnjqBg6pU+2j1WUEV5vTBRwC1A4V+yI5AYVskJiZHp3wTmU+BgBzwqsW
ynMR0UEvIn7v6HUtpkOdW4II5U6EX9HnxAYp/vvOmsD9pUc0BPW2RjTFNXfdU2w64yBk6634d+hI
8EgHDvmUpS8KTF+QJ5GHzfmtCe6tCsM2Af5sWn/Hf/g55/nWtWonRKpUFDuKMZVvPjCV6AhuiheX
UmasMGl4E5A1pNDJp7CGWkdCsf//zhF5fSLIY10ogBImfel8+XBoqKUStjYooY2MdLwIZHlE7HGc
/Asp29LRHcOwFeBPVuz6vnSBacvDVVm7lyQx8FTSFv9wjMInDXMl8PVI2OHZpu5T7b3xnEf3p6c9
EEalwybZJfbrFI/2pmsdO7pBdO5OPfsdkpgTO9JF/lKN9oB2itvARx1owx5fQsGbsXDTjq9vfo9a
VKhA1p9Er81DZAABFJhekIWnyyDozxfknAimvjWsM03Yp+S4K8x2lMxXN7MKUfvDFDOsRGkHzBnH
txieiZFkiZArK8gW/+YRaO9l0cZuB5mZmudJat3TshnfSWYZNF7NPLTkMK/LYayXRq8QJ8/2pjEw
IF4Sj/FryTvpqEVSqCWkjs29y6W3YI8m+ynkrn5yXLLEA57uLK9GBTouDP6NZyloNaa/R8LVZBPx
HnULtG9m8c5vHHPLmK29nc7vU97G+OdTKjWop9bLILAMppRfBqPNbeKg6zYzLQzX4Mtv2uiH3zd0
sHRbKTo9KL0waVuWS4kesl1GxiA2wSUCSNypJE0lRGKtdAU5eBcOXHERzC4GCvNdw86CslY2lmKA
qKA7OC1PhW9QbcYNxSn5pVT/KjaxoXwENNUhvZ/ZXMEX8R3Ll7HbyS4YC1KiZ/hGyWz3tPppKWMS
1MW7xqb3mznFEMdK5ducgEQ/wyFUeISusl42h1KeXe4cDNuvQIrm1gPAtM+kaaqR/UyNEf2LJKrP
ueYfqAj1PzLsizwjpWnm6PQn58wpUg7q3xVRRFpi/PlbR/revfZMhqtrAAmLK7KWo/Sii/+m48KN
RLEmoKO94BD9V6ugXh7ESEj8PiKPnRBaGH0IoonPqFpIYic7l847Mn4z9MubQ1uEqJAQQSdahiGk
zLp4g6Fe0kZ71Nfiq+NqbkoW6C76rYn1ZHBoMOWwCYGWbQjLZrE3Jh2X59PDWma6rQ8Cj/YSzoIP
vHxJl6WsXWA1OXLoYDkMOTZHwehgo0M6tw9HIMx9CyHHGUo9Sme44FJobCcqSdDU4Mdd1pxT3ddu
6QOCaSwVZ2FgW+87W2mWDZJ65Azmg2FDH48WpISt0rJ4K+yLgOPJMDfGhRwSlgPHsCqlclZyott1
0YI9E15kVl2ZFsu9Jd6IbVK+MX8OIb41vSDcRUlqRg8C6Ytdv5geLaCfzex+2x2OBjI+LayYV1Vy
nHOlj1RYY9d4ZMG5Lb3S9KXEleneOYlVO/hy0bPKBIiQnNSS6vCCtGcWLDeVvRpamn9SJrXsLCq1
kxZAYrP3g+dyzo6I4U0I1ULre70lp78opbzyC+WhzXEFW70to3n8YMdnZjjkBmNclTKWPCxWspoH
8iFofunZyd8DwYjW16JVz4L7mLbXdl4rHMxdsGbejpXkkqVYfKxhiUu9G2Fggh+vMuPfsWq/eENX
N7O/rrkCGQrrDJE3Jl9Odud/roOJm95Vx4JHx7QTt1jqgV1kvPYgMpcc63JTjf9oi54xwwyWEsg+
psVeYA3rQlg/qQS8HE5Avs3vrBt20zoVoTiQ+HzH3QrQoycym7b7ytYyLvltncXTtgvIId0Qlsff
co1QfiUw5iVGvejjFpQmCWXF31n90zijja7aigq9Eego1IVFqgNVO7R4sWvnM6qc24pikuhAhjCH
9vzzbDdQKt9rRHfNKso/ysomygliAXT4lpz/44qt7MSfn/2+PUKRvA6r5dGZaIp0tSr/gbWjd4Lc
0sMz9B3XBXFF3f4EBR9kizHu/sWD7BK333+L+Xw9/RhQZOKyhHhs6PCYr6LOl060H/mHXQ0nuEfN
Zs1ON8GmG2CoHpsLSchPjNhgqRJQQc0Hy1DZSGCkFBfthLQ4DwqfzIHjFKEWOhwh6XJecs9mbNaF
uGcHZQpQ0Cltq9mftQ8d4oF7Tmb0wFJTSQBpLtiL94Q6SGwnBs0n5MQZHyY6T9121/wa7mzu/ZBb
MInbLOWXoCl9kZQTrcUsYr1ZNufkuDxC0QGFCJj251G9zlpZi9S5oj4ZlKg7Dk/Oqj8zYzIuC3ja
KnKG7H7x4PrH54RUzDBQOalFxzAD5s5WebXj8KGuxj+BbN/RKSGfv/bvDH4AOMI8VPu77LhDQF6f
8qlMlIyl1RJVuqSIo/facfnLBYgwZomTmRIaBhw7FgqtEVifJJ7VPURIU9vpq7Wk96hmEJy3Moh9
rxYgYQciBN+84RrP4mXhCvbHwQjKUFhMXW0AmwN1N4+tbgPSCxaPiYsUb6lp33/dDvxONR5EAJ81
eM6TJCc8vkb47gkVsK9pWn/qaJaGDrtLxsT4CmbULEeEx8PMJNi2OIosmKI5NPvU26LOVPDnG71B
9mXf+7+jbtudJEXzLsRgN/zX0oo+G9Mm9+guM/DYpZ7PyZiJTJKNP9jdluAZM4Sb3wUXPHdljtpd
h68vQGR/PZq2fljyI9jMKqGF8K9zORZ9/m7qxxLUNpdDbnFhb2DEXbW+swLUBWdf5SQiOG+gNxne
mh6Q+gP6E5m3Z9BNAuxPVofb97rgsKObJRc+mbjgrFFGW4DaTeKQODMh0YRaR+hVJ2opa7rXWbV/
sGXF+yqhwwwSk2fR3IqV+65bvB24gzm0d460D5od9cSm5v3UeChUtwurtttYIIM1KCC5xnGG33nd
lJfEpG+yJaPdrW5WiMi84aIrMcgeUN0SAfTNkI2wYKX8Qk3Mj1YCm5bm+HHPrFlpj9zMGmSVPspD
MA+x42AkRWIL3eQyfHkNaYILoZ6dUcw/FNfc3AZRei6cHWGezDSpaNlDOCb4hDPQHuiAQDK6JXUc
XBfYxdpVcaHpLL5EcN7bYhzVjbNgwXYcq0CIG+MaYNpUfbrbCAjMR6CM6nDpQwsqRd6G5Q+hE5nm
Jdl6GPHQfMtCHT7P2iAFjta6Wrp7OKJBqiBJhzk7HgasV3PYFtOvuUavRK3sm9Y1hshoifyRg7cv
G4MmsUj3BGSBnJxJ79cvHx+duIDzuMxjKkzzbgLQytpsgiSmMklu0Nt1FbCN+w8ZVymyqD0d4JG5
/cNHw46c5Q4FjLgXFWMru7sCx3ew5YxyE5W7YTq9R1lTGzJmpAur0HBt/GG7g+kkEM7k4moS5T7p
deQf6fXEwfTczdndJGu0oiLlhodk4eZUTUsylAKCSljrrBnVO4eU4H13Fs9X7yPJ5/5KeailRnB1
oOk4RnUK8QMHdW6Z1hl2yVgCUjPIeEJ62SWfbELm3aKH5fpgswF4oBw/B03KDEEgHNIVx8J9miYz
ZEDxXLVYl4F8gewqyCrIAa7VaS+FkTr+EMZQC/g+sBl/YzSx9OcK6C/Ap+KVxGScJm75RUXGy0gd
ODRmZFU04yA6qBv0/ZdbXq4JwG3NVYB0ow3imlI194VcmO6mLYvhGS0zLDJLSEhuaToucrgjrbu7
O4KjNkUX3I4++lvQjtoYg1nlX18In0pySFfAXF92GNjDXC7SVIv35XecygVtioIZ55oCEdYTv6Cg
xH25F4N1e16K0vAD1BiEBpi0YtEl7Q7GOeeMUhc6p7ROi0T5OinBRvE6K0NR25eRvdOol0SDjcME
fcEiA/WKTQFs8GiTAOrnQkDvpZ05mijqUemXIu3kXsTxvaOKeZjrxAgihZg3BnBhTdaGKIhQaS9Z
quKtCQS7t5apio/baulvL9m7XzFIhJpxn5Vz2B+yiqol1onzLh/0PveVlPiSg5xCm+68AW7ElbDH
lQ9UJXutCDvDcQkatyrZ9z4PemrYhGFe5hTgYYTN3vqP+weyEVGUYbrwiYUuCgMS2qL9N3wWFTKl
xfd1DE0WbRCj9sd9zi/IN6UKY0olw0/RjzovKu48QrbkITmCcHA1ztXjDcvX29MEL5K9/v882Nlm
kJjIKaUH/fKZmh7yOZhxrPXQX5Cjq2REb+DzARxbwS/dBVJPXvpy0HzZ86j/7v794Xu/2Ksitr/A
rU63VK9qOMXGNWmzokNiocAG20nwSIeKxToXygooiYMV9QX0vxzTDp3TNNmUTx9JpTQRq73cEEPL
icRnatbciRG/Y8+1w/MaeVs0as0xcZZRDMN1knZXk5qCgE4LMr6tzh/Da8plC/BkZ9i2ISVHtgQ8
wdRmfVjbyBbKxPsW/7nFJCLpKeaOWaeKwbu4whxoRE3cxNwXnoZ3dQ5q65KHFLdWNHgJtC3sajMq
5aLhl2P6kwwCxwUUZwFe1Wd5BUl0Nz8vmj8KcFaU7XOnrUafIYixW8rbL8VTcIMQEoM7LRWiMkJB
Ve9RnAt4kx5iiNhE2iAIioPN4Be1U0D9ynWEeo6B2qYXt7wt0UOQamXsy/Z+Uhg6w7NarVGHGPsj
5BLdh0qtFzB5u16wjVxPIxIvRHNfatxOpYHg600M9khFR+nl2gPsG6dXGUXtsjkv/uPDIhbhZkFJ
Ll3HIhK8ox242nSFZHRZY7MPU+JFWq0ozuveUHdFkQYUoGY1qZOJpGUqazPbiWgy0JiNdb4Re+Fk
sUrQbp66V15ZrELb5jsylfgWUhFD5JZbOGiF0RP1spCboxTJQ4PcozOsDtdOy9X9C3BI5A8V2H61
tZ5DNNOzePxEbUmko2tBxUH2udIhlCnRp77GnQkhwYcsBHIv042BIdfnPt3CmI0HPha38SxHCDjT
cLs78PbYx58uR+GL5kau8B87THbq6WD99cqS3ma9SbEKaLrZIgaJ/1qZWq7B4l5EbP5BDA2+OWFJ
Ne84aUqto0NUquGQEHtsRH2Jin49+t9KX9EFJ5d/XvG3bGbeXJOTIK4PFxQNHvO5XqsNUkLi6vLJ
8FrjrS98/tn6xzsCWKD3mJEWVUYdxwN4FFKR1x7hrdAJA09z5uEfWse0BfilbHXjLdj/I4Uls7gp
nvb+MhOK6unX8p4n9qoR/DKnBLSGOOe/jJ3xv4OCtAXFp5mH09haltbdfrfgWACA3A/Wtlyc1CSj
53wNStnWDdvHVnJaimmsQs7aYYYZgR7/fcQ7tYBbN0NJPevPUu246TlBADDS7JVt89CcB4trwqU9
5VWdNM3WKpjW5tEDhevU4UFuKAoSQUOEE8tazbg8GreBHaRpXHJF/g8FamZXjKglsohp5Zx9PXRd
UB0dcHxYcgQ6xWUgER2AzfZ6BBC2csuhsRk02Y4lsVmqpngpLevzxFINTKrGVUrFVsFOa9QVkJEc
QmTlV/0MX5IVXZDINpfgoHDdCZCooop23GdTnJfMFBEcYmnaRnl2vSYRI29G1WkaLugAXRyQtFmE
4sCgVb/8ORpqStuLCoK+T7do585PtkTiPVRCY0p0S67mEzKekPo713QhQBZQTMx85YVsZZ/x2r7L
4nAFzqKjXLqzH63IicbHFJGQAylhQjmk3jfYnwJ1497vS/AlaL77BPbYjfez9TB+pCOnMSDqKbWc
uIsYckuU71bEB7mw4zWc/xpNyeJl05/wjoMVC8/bQOVVgljCEJa4EElvchjSSOjWJEfMTsvSUbdC
8hcWTM8AMfbjJxbyS+zPNxXuIJs98rn69KQfD1HeXrXIqzgDZpF9mB/DXYQHL5d/Z/jKigp5fGfx
hALbtI2MVBaxW6JJSu9oHcLHbot20ede9iU4xLC6KsL+nHWKDEJbDO5ftqncuGE86u38lOjg18Za
YQLtfncgRjjlBd2kq1hDgzBpze+K/P/YsCeJmyOTSjWlqmbUUObz4NYp0Ic3WUD0+FB9z6ou8Bht
2fauZBLUsNELNlw+aALZ73PyC8Tme1sJcPdkpB3tlJXRw1aTaKOsqjhtV0dtNuS1PbdKaGVgeKGX
ICzNqKRVKqzK+yRvUiAu8tS8iZU+UZLK1Cdc/RvW2Vwi3g2G/gCUHNilrcCASZhc1fItnEbTUXdo
uM4cJGENh/mDJPhK1A4PBNZxxtaKXU+WuJeg3EphGzph7R26VUJrIr0QoF4PNwtfxWyx/bpbdPOI
RQg1gFNmbm34qcW5F0xD8U+WTEaex0D2VN5p5SmlQpEeRTd/quMLLsSXNO6ik+Y6PAvg4xEnFMXe
IjDrClTWoXFxel/3G5GuUK45U85O19q1IIBfg5GT14LNmqfbpcaxVqAUOp79XRJ8RhWu+EcipX1g
crNCLri4gGzbQNZtvCw2g6gkvWecVCPjKw9VqU8YG60VSqiJ0aLcHPWQoZtW6oZzPzgTzQrTLYCZ
2aMohlDoxRDReh/y0xGwg39/l8O3pFWxBv5oH4MnzElTKTd5O8eRskl8F+9pu6kRLIpWn6AfCyCj
ld+nhJ1Obk8XpH0gu9hJAPpsVNH7cFrBMfWJyluV1Z9LwgVPu7CaAUXrNr3ccDsEQhPyL5ekA/7p
aO+9iCvz0uy4LDGf5zM5cPaFGs9at5XraFC7VzqCGvUz/27a/jpxTG7PlFgZb2Q3YMzE6pxBOVLM
e6cL9/Z+IYcNg2pAT/wm/tiSq2wBr/55pTt04bnCACNaFTSWeYW6zjlT7dgGNzncKjitdhCYFpIO
3mmHwb99BbWgj0YoIrBPCQK3lvVQ3AnKakigO4WDTzU/+KkoQBHF9+H1i8a6jR/r8Z0V+VM++02q
XrP6jCPdOd9R9gBGd+cjgUskmIfzQU5RrdCybh5EwGxgq42zrLh+94eVtYU1Go/O82TqfLP9UrGU
fiRBIzhy8+WAm+7suo43x4dOwstEcpTURfdXN+PzM/lyNXdZgfsHUcEl9x0I39gwiHvjmw/+W5Ia
L7Db2dEW4/ssMKxcfinVEk5Tz76f5EuwfN5olU4GNYkA/UuKSblXs7+g35cc5cy1QDVRkxaWQ7H9
PqQgs60itV+7osmGGRAhV6yujdwyK1clY42PL9ttcjXB6b6IW0sSJr1G7UrP3Nmik7duM7Ryyfex
TLW1OOQMxxtF8vOzURhB8Hl8l3Z6D4iusMPvRR9b4xLtk5R9TNePBgIjyVxhK9Rddle2y9zyr9tm
qkDlL7SxjCHy9rr9kdSu8IWUF0I7IjytTx/s2edvRDGI76244bQXfnlyPNhYyBmTDWwU8iOp0Upr
hwG0m9lMokLlQgx/B3175xTTxkZoaJtnzh4+hIulFxPufIJWd6EkhcwOVK37o163FOZYglka7axz
O3R0cjy3raZ9vxgIW0wrWGKnwSP2szY4kyPortQE0+Y/gG1buM7xXN0XzbTIt4UUEXDSUiwGWAN2
oAwwi6WxdR3esU50xErhKnDMMHC2xYE/UqBkDbIl18kJYeoQitHtT0jMn7122y2OB5itaVxUBQbq
oDBiAyDwpG2pgfmDoqJsHI8SotnFjQkUT3/yMTjgtai2msN1ZGDty0igHA73ITrAyCuzpou8DZTx
neIakM427T6PPBXeR1LRPRywzi5jbLUVk3lacn2kCLqh6qusdLid8aXDvVAErux/PtYr+apT6ekr
BIgXdP5qQdlvK0/vx62g4VPetI67/4ytDIncnKbgYVdws/7QnP46y+plIANbHAaBiFgj/EMPe7EX
BzrXk1AenIxisdHfh0k4z+7QGPxmzDESSbAA2Aok6VQ4tF6GaKtYmOmfHRKkfWgVwZdm6v2AJCjl
Cd7NCoadsw3ocXjPui+yFxAiiPkqpmBhJtCJxTo48kkxxyjiK1cXSvgEcKxZ48sG4Wk/UJzr+6kM
o4QUUQ7Utp97EpeBes1o7Mlfv2jfCScckFfkCJ0xMzn8yRCJ3KqJhPp2eXyoIGGdalWgb+DxxxsN
o7QSw0Xw54QNt6d1KAQTyfDfNLa6eoXFF+IkeN53NK4jkU3YOJmV0LzJCVnSK03CNjxPj5TlS9pG
gch1E5sCa6PM6MVWoGEI/63L77t5SelJiDk2EQq9EmOLdcKPU5Hy/4IHiP8JeDYs7kIxJP0qDe4x
pULvBB/W2jbIo4fNbfk9Sa7aFQ0/B/jBm1tShpZwz6PZH0H4F3k9VT5UHgFMvyMULoe6HAWM/OQd
8ZLxGAMd0gLLqSgS8LR1MG2OWrQQ3RHamP62tg1BVhxgvy+c46xhhAihZVk/E0c3OTstiFDwmI/W
rHbFDaA+I9XNvi7m57g+ZGYClRMJY1bxirWXcXcERN3UjJYy+HqVhcIt0K5gwWu0gQrpIbf9OShp
45ZFdBQfqR1KKTwfJEdItntLCgz1VYgot+Hd1SJnloiBEhJ6EwWZGhn7L9Nz62dk4cn9ja1cQnLl
fzcJO08/wnHpJOdfIYomsD9eQdG4bg/ZdNoxKjMXhitkZYvekN5TkqDF0SDAZYqzNwmap5NpCoV9
m/eO2DUGJfRtfQVudQkKJUh+nKtBV18H8IJSnSVJaqSYXyG+lrvFkAX+o8LDvcNQRrQUJGys5/GT
44m3ux7Sa4ePhg44PAuUqaiOhLc6fCudWpV+CT110HxMsLZM2cQu/L3cqvSSa7AQvlSIJTC2/ivA
o+ZlU3r3uEWM9goG1jrKzXKY23znIIulGL3ys14Qi5E6fnicDpfnisXdC5sLQNVHVDruivvS5z03
pjtVl6SeK1iMmHVZuO2toyRTeVh7gNi/dqxOeW0g0GLcZXB5UrvpQIbnCyMTU1EnXrJC+uMap9u2
/ft7ZQH8WSlcjQaG0al4VI1nW8sMlAyH44AUaMGbK44bY+p+G+bsyqcA6dhUtvvkVdE23TZUcTl4
FwjjDaiSt9ZiB5Jpspv0iAD+gStzODXku4cz22ErFBPyIamJ8f/ZaSu7HrZ1rdfRRiCV5CHeW/bM
3J74DHNACsKlLh4NSYXEhnGVAEmCXyh40EeAC+Xw5CP84XJ65ctJbsmWOnsPPdM5oBs5ApcrOtoY
6PYd5PxWIzRGxxKfureO2EoKcrXVC9E+vvGIRAeHa6W1aYpxwCon8eV9REiWmjRCxhRWg9SHMfGi
FCTZC/Wog2FrPpm3jDeJXBoG9NeZtgBpJ7CbLUbGoKdxOT8lErAf11BjasPFiCD7a3h3F+pQ3HPM
En5FcatV4/CMKtLkvOBtGnvGfZN1rkXmz7PJAJRpGhtRHt4dVNlNbggT6c5SPV2FII4xS3DoNKH6
QXutzmOO/TBgCeUYEE7wYcVHx4bgkhsry18julq1ywKU93kOVxDsUBXhJolopdpk47AQ9FwR1he5
NuwHP7wwgKo1sOWc1oz83o1Jt69X05+E0dOcWm66LYSkycG69HtBckbgToxXkfFQGW4EPNk+tjUL
fKRuagOB+pslPuDMHWiSjpE3cWKjnPh1l00ZIycuJaq+kLLVhV2VghMUTV8piB4H1e4+qv7uve8C
91++0hKLE4pumExTTtKoftxDHgNTJ+Wcp9JIqAXWBV9oZ9c4GY3QhOgiI6BD41n0jhH0wSSVtl4u
dF9jh0DJxCQtkWUnCSyJPXCs0O7U6tMZquzgZd0O+Z/g8/9IzxD02lh/R4btalDyyTirLF6qNnhb
5VPp3dcmvzEGT5r5ZQRINgHJx4Dv/1zpONqe1FC2C4HeNm3zq23gWEUi1Q36I4XRet+ATMCRdzRS
2WhrIirGXqGcmuYIzB1F7PxrmXHcaohLz4DXF/UlYv1I4iXAAkVLVVfokDoK8Byrs4c8swOGUGv6
RbNXBTo6ZMlRlYRRGLw/brT78N2ANO1i/lyGi1nUPiz+6Xidv8nkuFU7jB9Jz2vZvOWWgOFbK1z9
+n8Ys4dYv0pu/fsFDQGL6p1dkqBjpPqCXCM0OoWJGw32wRdfnjo1mfojD5HdupOcvUTsuu5bDviv
PYw5PQc/QLkikmV3g1KaUmh+DBQNfbGS9R71dTmhgGmv48L54LuwZUSfmpntJ2K4WY0cdLYx0+uY
PhMKh5ZdPtT/lkkUN2SklhntB4CJFn91RpBdqueUnFWkKSBvbUK8eordp+EOzuuGy2+qMF1C39zf
46mkN+BauQKr2CDZYzTKaNy45FxjTdw2R2D6s/qYgnkx1LhQanIYgTsl20u7AQu78Y1PmZRYhbRN
IUZm5A+ihnyhxLDrjwm4oh4IZfvSoqxmWgq8IFuDUhj/JjnE4ZAO8BhDv8qn7AIYvTKWgxlJMGBv
faYTXzfAAq+/LmDbKwLiuM+C21Vya2uc8R7uJuU6Rv05BJEOmQnSaHf+K6RsjQkE6QoC2QNdHz6v
H00Mw4QEcfNK7Xo6WzZpQSLMNGegKO9pefNmBwqfn6u4E8/K0+7Vnfn9uHXLKVHbtpgxEyN3CV4O
mriORUgLAGtB1W/3rYx0qOwDdx7/NdQSikSLD5NPk1+8pDNdEu01aTmMqyjhD6/GA9KGvuZWlmqT
9RGSznLOFTT7gedfku1+nmO2T6dNk3jghzxR4oIn6nA7QPjoQc+K4MlUABm73Qaa2//OoZIO4Yk1
Lg5mDrAVUxBWqJYlFHIc0XG2e4rR5p8qBy1XSeHRX88yXN0DkSe3EcrjMalEuOJLa2pHrPVgqOY9
+gY5zMtHahgRk44utwnJLZubc1DwS3oDpLgTkRZ3p7qYm2JpxAyzUhFseQyTKOZ507jFFXvp8J2E
4ea4qgAHIhrEfTfQwTj/i2YhLyjZwmeUIdY3PPmAZH+mTLQ/arbHOxe+UdosMIqYSsqACy/ZocbO
jIQZR8REM5gpJ1ROEKdEKmXzDXEH2AfSgtPTxF9tRGkgVOy/huEieoqRHdoPEX9aAZAvewsHdKC6
weOXPtETUB83ODEmt9+BUz1cgzOtoY4qZP4xz5xMhVDQZkA61yaPTrFAjskvUmTk2nj64ZybyDrw
GsNtwpWbQhS/YmN4X5UfkkgAGWdWYOcnugi/D30hWn4fY+P31kOmNoMMHXTjuUWeqLDZxxekouwf
CnBqaW0emvEJakD/4xNICsE7ZVx84ZZ9fALbtCfpc5OZjjQUbItI0bdo1iVi6pXAhg0CLdcxKpij
odUAKwOG66Cb4dTRtGkKmT+UnSEDdPzgzISWPJUCDDd0hIghm2LSKzEkRI0CLV3FCOKnwUqVU6m6
I3vqvknFSb+VSJ29HP7on05bA894A0WDDjXNCskfRvagZZGaUI/WuOtMOdibxoxrUr4ED8/vQx9e
tBmxjHIzWR6b2R1VSKwRkbt9TPnGOD4wxLlsX5PrqeyjTG0nXC2PiLPuzXox+yDCUBnKpIxUCpOg
2wX3mK24eNT2Nk4IjBL1x+mhZD/V3IOWlNdKqqSiI/TpuMjGS6U3Bl9FA6YTyxdlNK6IRkXp5SUT
qjgF8wZXtWbtHYbvSftBPm5J8KiDoUO4ot3k1HE/i0MZymdI6GYhXOIVyHYC/oacFR7Ir6s4lk+p
aD5u3UkvvcIYWtcMZAH+WoWP0ltggPkxtm35Q+4U832NUiJTuQKFplvXABvrt5/O7ztomviw4neA
s25GXj1n0o9+RA/kZysCUfBSe4Uf3HGdbY2Syze5Kdjot4OU6I6xBII3aHKkDSfx39GgUbgsvBuw
KH5f15LpzE6DEdtf59FHnyCh4YWNL0Png+gefXf6g8JiNCyWBAISMFm3GbJK3IpvEvod++QRk3Ae
oD81Qp3/ROj8DTw65hRLrpGqChlHk8ZoFES7ri5TTgLjNS2Yj7lkgmRybSGWE4GKLjVoUOuDLtJW
nJ6M9BqFHfDRiyeWKkUV/5aVbLhL1vEF9twPGGr8fWCxBpIi5NvfE8WC7YuefPEahzOBcc62xVJw
8FfFQLZEgVadXFOwl3A4tqJy31fwx700mphw6HeTvh6kAfCmZ6O5MN+asFjWwO6liq5nagzNA1WN
5ljk1Y3Iz7euCwiYsPxPHlWn0snYYv5DGo6WGo15wiKGWcWyiXCUNjsMf01j4/LaHAgXjB9UfMoR
1F3fvMmcq4SWNQ2tRZsIs4NN6xwRlkH+4Ue36ddfNaCkxedD+lt7jvfJxvJBgiPAOCDIzs15/AUH
Fj87zZ7VQ7ku+/60JzEQFnXngYGkUIOUq3B9DAc15vo4vjicb3fgLLv3lLqSLQAkI3+fvgFLkJ+b
Js1KxaW0m90dErlfzG65Xb7fCebhxeffox2BD7sUmWkLq8UYyURgnFSYhfh0P6bsVJEyU3cAba5H
eM5yPjR9G1Ct1/tdiPGXzgVv2a9UcG3CvExAwE9LV+5wtubbIvEG91RSSs/QcGg7JpDGeG/z2rVP
L3vOVqWfb2lW1BHCPD21RzzaydM5mUMjm2b1h4hu2THuCSTQO4m2wzVxGBN0ty+hMuAKO9P1rwsn
8YVs36Rt4bNVtjQ/DHQ9a0uk6ffVunl+iT1yikz0o2PIZgXjktHW6oAmH1oc+o88zhfNB0srvUwQ
W2O0FwpdUsjeZueNmwErcuZKX308tkv1FG+HPLRJr04uoiemyUe6h1uvTUqwleOa9BVSDcHexnpu
O3bYUsHLUatn4k7h1lP9ExV29hdxUdkATYF1dpY3Rz43WOoSisQ5n7GlZyJE9Xw6nZWYH2ucTy+P
dgVA4/TlenDw8/0qWQuHBudJBZopjMI5kLZezvCS3guSzyHgQKTQSd+YwrlHreP1iZ/ppwr3RTW4
iVpGqfVVyepqiJgwVH6fg95heTUO8k7PmIVa/6vTqM7Wxco/O/18KYn64QcpRXSUJWN8yzEVVWRR
aUWraZefXkjXAhdnRkWIhPnwRJ5xjdG0us45oCujHzgLsyGNNERKPzi5CkXA3EVBonqrxLa/qUkG
0f1IXih+bRJiqNwaEGiQTvT4tk7f9owinjS6cyy4gLHXSUqbQ9KitonAH8EHWXcE3pcuVIMmWaTP
z0LbYjztzN7OmGIIia6abOy+sbynx13yn95YjhSKpccpM6N2L+hqMPBruogVhhBjBB8fSxP5QGRh
hVdK6eeqb/hXmnppIUns+oe2a+p6prQGNl+fbXcro0zkV/pA3oxxPNLR23/U8ooj5oiHoRFq9+L4
ZfyCjsZmIR+mvMZR9NEDklwPdPlwgvhS9smnvKHsBcWwCR612wPC7aqkKH9uy1O5PDtIQAarX523
B5Ry4c5i9P7I+7A6XuMx53Degpg6WovS5b257SqCc8k6VlpgdSBAS9cPGZ6eJONPlycmU8cmxFdl
vL0VhTxZoD6S2ef/xdZe4iNW2sBDudqtapGn+5InJnPqAtcYJ39lcbJRkCCBgt53zUXQTGFdKZDS
eezcsFV/XjcdipoCdL1rbrAX9RaQ8bzRIq6jmFYAudvC6GdpyL5IpMvL5+RiCsbMY5MqyUU+THuc
ukEBIJQA4cXZSG9vET78S/eakOiUk+Pbp4PMut0CTHMvskDE44wNK+yukgf3paP+Jkc7mIoyBeoE
qgw2zH2Xm/6Ec72LXn4jsxzm1u/sbyYzU0h4X7iXYiFKYfucHIx/JT1rhKL2P3sNdfu++kV+kKxe
Xy1n6cvMawyCSJE7mLi/NEWTXhRi3X7D77hePq5kD6ki2ZVtsw5aEtiTNyjdKDo1dlX52gDEHyN2
ahObM6y5GrSeVS5XmjomJZu92rJWoSiFhchm1xD3wjMUrX6rElZwCdsY2t+kiHrqIoi6wCi6DIQ3
pk/FmsiJSaJU+GT/mzrAdLKo1pilWWTA+P29OmQUk/C9GZ68OTQy+XJbmInsQa/aWBIJ5ICS89Yf
QBDwTeTnvk+AVTz2cLHu5MI1+bc4VJLDvEZemx0IKM2kIZgBwPetwR3//eGgnVG2RXm7153ZqVGR
15zrieBp0OjpeIiwPC15wUl2sYeNtTvxrjYVV5X0iBO2Ee1nSROrEcUzEkLIMwnlqkqdwnI0Dt0i
dU0aWYO3SfCsiiGaTII/MDext2AJm77f9rierNdun4Bn3whvVwSpUoByuw1Eytlcmr4jk3eb63cq
6gpObGqLOb8odBBzHTE3E/0s/DLFAcy0HNY0bRpIFfWawgHVWxiH5sow/+ePhjxhTdW7ZToJF2r3
VfY0wHSgY1Tgl6c6Hx8dP0grRoG/10YAXntY9OsZWANRDD+dtBSaecbGOqcfwH1BCu7NVP9/giI8
AHma+Xk/LjlbZ804yVpb2jPVw8DbTK4PX8V7dVUROJggyX8p4130hNmFilm/VsJkqwH42o0ZH3Vu
SQzWGHZ2lBrfCLdIVq3x2T1FX+StZW0gRHsGaQ3y9hQwnRn0T110Qzqbnxrn+cwE2ngDUOKDC5up
hzHeNsvnHoYmo5lqsw8teciZzBiIzD4nvHsm9WQ1oJHF3bASRA6kQH2Q4m0IAJgDRRZwn8xRGe0B
LwpLXkvZ+l8A6+p1us/QgH6pTtY18GWj/cnyhaYv+q1O1BXF7eJcYn8kbIENCuwqQnnbNcRWN5CP
E2ro0MlR8gy6OWeQqg0kElN+0N4chdGHB06QPOo1WWCC6qI4i21LBKPrjD1/Dibt0zjYZM1+plTE
M38xVLobEIZYnZrtnmhkvfumrjZ4vX81AzbcmxNYtYkLZpQ+9OUR4Dl1DqninC8qF6ngc496NQW2
EZnLS+voMzZRWxyRuoLFOTXboqgO05QwM7chmwVWaRtxwCbJXxWMuNGl2gJ8HDm5nGk7axs8qTam
AL3vOeYAht5r0iQOpkMVlv991I+EQB1rDBFcecakyX0y0FBhydIWogsjhSrBuOvcCUxNbxcDz7np
VGwPoaotA8Sn/RJoPe1QSsU/UO181csC/UJzhswAH4EDf825k/vFtQNq84WD7nVSZ0ayg8I3x5ap
Py4cIEgRqNGrbaDiGXMuOzrcj+xqacTqzYok0pwRvk6UXcWfy7pPprKVjnwjYMylO3MuygFII8Z6
oYBJ7RtOZWTl+FrgdnnIuzXKQBcQXkLIZ2fAr4DmHq+1xLo7IVBuHEwshdqY5/fN6L5qrnNh+Kvo
oWamh5UERDcKduEux3icoXY0Rk4a1y8kzHXG4Plws6u/nMQaPtlBJhnICesjPjJxIJHZ24QOMdln
S+WbftZHKD0Hatef1KpKn+U2YpOHce6twC6CSKv61C4eQNBpXQf/1WhbsZI2hbzY3/eXOyjpzpfy
PTL9XqFQTTpXJRsAFe9WpvMQmTjZyhbSasBfCL1nF1mOigGGvPHGcKmdpBLNTRbNJyMJKV6fW2bX
CPSxCVeoxR2/WoqZUWhLezdXQb/okCHVOCs63XPMJN87VeE/SrVJmzg5eqtqg8y7pitZKgr+hVna
epjGBBvSNwPotCP1Mz4jxvgsqFTeHIlOI8QRi3cJpn8/1PVUOug1KKE6bUPkulUhBs6Kqs5GRFZ8
LwO7fXOSAVS5bq7hXmjKtDR9sstiFVqn80IVNAAsWz/5FVLNiwGy6Pw/LLtOCjIhl9U6bxaocDAP
WgUODUM3RlS40thhyMDOXR/f/kF0DI8JSeBlykVAc/IkIRVTHa+GHBZxq7G+hvU9bbdXReAlUlxs
HPCJ+ll8wUOxRc4TxUqKf3x0lehH/9w7gcCmEhI+D0nZyQ+OVfzCrf9pfZE8QF+hywSaenQ5ycoS
EionphqV5vmFaV+hYeLye2Tx1k155H4tTUhaDgsFomGVKGDAiv4cQci5YKJLZdW6+tcxn1jWcyA5
dFDu/ptcMIepHOC8LrbmH0Y7PyX5ljO6idESXh79OlFuDfLwKdjcB3jQMFz1mvcHhZ9Aafr42wlZ
12wj+47wiqOZ3t0Lrklf8pnH8Zy0+pO40SrbpdjbDZLiTTx6Cfys3ka3hRq7yC49DhHUTzTYDo0W
E5tTMJiT7LuBcqLoKzy1ds+dtPFzflOGsAREZonpNpnNtpBIRMgSswqwVarJUQULDFaBIuWpCBVV
KhhYqPt5X+NN/aaFBaZxudWxTyOXklWYgWazxQ26nxb0W2+q09w6I5cNVcBBcH2BL8s3VD01ARfV
Swf29PN0HsqHeD62tqr3oEwdwQdQTw8Yc82oX5LbWKmtIQwM/m4ruf7v9g0uUXWt1nm1D9vmRDFQ
aW20FcN7qLLGd0VlQ55P5JVNc9F1uW+DNBIpXp5v5Emss3mvnZbm5e5MdC0q95O+1rXUE4YOHYcU
4v2WAmZsX2uxMtbKut/oxa1+BQ3FBHynjrCnRcV5hzpSEwMYNrbnOdPvhMxQ4uYr+I4JuA4NTl4V
IUIZxIO8+noXvbTdEoF1J9vWg5S7Kfwve0WsP/5Zbt6psUfd2APfWpJXUUT4Hrh9Ksyx85hnfhly
P6PZC5h97ITvM4EufGuLd0uQHhbwK/Zal6WDMu7DP65DX9qlw9BrQppDIi2pCwp7KS/CfYeNlbnO
Ylh0AIHykRpYvAVJe5Jcz9V8KcfHpqQ0nmCT73/7AhoNzZFcxE/4KFFSR4lx0bpmXE43K3xEvv1d
6sqsBheKSvxJ9hNdMaX58kKHKGMnRpDEw8wvKSVp6eZSJMtpAs/fFYIkgHEEUFyAj60qv++T5/v0
fI13G3iKofT7m3/bHrvwDoCIvp2LUPUsFRDq/YR1d/oq2lObg1VB5cPt61XKhsmYnEzs565ap7mX
tkHkx+va7tIwxSnpZmwfoO/swBEthKfHjG9dpTom+35ZnrW8UppFckvqL68e7tBy4sO7QQA9Zks6
o5ifd3gtDNhI+4in13fWg1lYo6O4DDvz8Wv49mKmIAJQOIO2rg/XypgmLxTJouuRV92c9pX+t1pY
Y5hx4KUb7nw4DOkp6/gMZEqGHwcbw1apYd2B3o81EXY7URJt2Yhi+1aU8ojeIgxh/M6C60iIpPE/
cwjauD7RKCx7aMDUjir6PqLfbiBioLuEwUXPMnTcc3VWCJQAnUGefddzvZet1qOgrpPPxw4Vouw8
jorfr9liO1QgqqN5hU4/eBbCIF/bWxf2/oNVh6ZZZppgcGfR09ANquVic3wzBQTZ+Txkjne6XzWz
JekhRdclmQ7/rR4ujvJvGfO3TnlSgsRW0RMVDkpT5TWSs975F4oeRr9bnsJuISjfnKZ98SBioP0M
VBimoGmvzHgI0l2ieq2LSzMQrGx5n/jdfhvl7BNHKPWnn5vVCWpTaKFYvkiv/SDyr3ak4569X/RG
MLOI2w9giRfIw32Na+XWvRyAv3HCTO4fHHFjIF9BsU7JBPeZDhpCq+mjWz01oVmeala864kYN6ey
nY3Ara6TvcfZAMQr6dtZnsWCAho1xX5HODXinHjZa3nmeUnpQNK8gtcyfFcWl4YeMJu9NWCNNlLf
SllBAG4gEOvWv4C4gNT2pupKzQj1BAPtrnt1KoD6B8lCFV270A0/Ux7T00pgxAOGpz3rREyMoxzR
4LL59fvqM86vT6JOmMDt02OtmY35W8kDFSklWEJy6NN09vFgRRj/WZZkgrYFvJaeLHoAU2pUJ8HQ
h8F7XOhBQ+XlkHpbWtXjz1mQ3OEAQ/47sInpi0kzjj8zbvdwjNLnoY7HWpo+8CpBD9a1fPaN0sYc
gmk9ps0EOzmz1mUr1zYTrbiKgdkLBIuvWlTKYQS/PcP9LB83BBh5Y/nU5vbVBulf1BJXomLPsiqN
+k3UC3YYpOT9JCd7fCdwxi1rbTgd+rXts8xa/vtXjN0y6IrPMkvp45cGhuuLUTzPBtVZawwoXSKY
2Tf6Hffn6wSUBWFB/nWRQ8kUBwvsmfw3Q/JnDt/m/TAvIKZfpTRRK5nsSQl+oobuctdwDI1iYm3L
T2Ns5frAGheqyJClzvJ5sJZ77XNoRNra0ic2P1LxqURsZ7W1Ns5rLwX67FhxHzS56t66Mc5JW/vD
FLHmsZ+wQaeiZY4seRbwz4tPkLTlUsZST5XRGKLtNeySMCpLPS9P1FEegfLcZkd6j25mKlpwMI/A
kHqhpQX9QIuS9YmMdncv1RUgvQzJp1NhGbKrjtFSN7aLTsYl+ZwBR3D26dERGeuqMX5nAAylyJOi
5jYNRGZoXtRe+CcXtMlpKZlJ+uRoyC6SxL4EpAMwbhjAFYPC8gfQyWupTNXyCpd9QbbfIWAZkQRz
nt6OGRfMEnTgcLel9w0pUytfeMnRY0GSZbKiT1eJN7IDK/GTcvHAnHCET4IORsc/ac8+p3kM0S49
saDQrQndLuuY/6t3iLqlGUdowhZi/f1LRLpcz7qPlaPd1wupLeZmndYQMbfVTu3EIf2aUmVbeMFA
cZW1bxPtnCUvA+0+06Y/3tXC2VliGVZtz6lSeQjPoAHpjaaA1ynGnkzVuhJ0SLoYD+Gp/mLeZGRi
UdiSiwAnG9u4co07AaB8SlDRm3mP0sv2D3cbuSnB6d0cjdnZ31p234pfQkACheuCTRNF36+FdHFd
y25dyygMLUPo2iD7Qh2Su4ZLmcBRwnNUnyDTCFdnHgglAuuJo7nbKxkcBZMpxrunx5RSe0NU6rxe
Ca65sKVNllDqWY89556MJxbBpYoCkMv7y1wbhiPGpYGKKl0X9Jd8y1l2GOed8Qv7et7JTRQr/jbd
R44nAfwkOsQj9AIpePbEkWQT50Bg6pIuGahc1Be2xUdQWK395/XepuXSKh6X7SiX+qUIqCUC9+tW
W36p4h4LuYmD1IvuTn15ePCulmxjCE5iQpYwopgGFrxdhat7jXaTPcpc+aM+56aQLGgFJGkXSCbr
HE0q5O1uVQnZLQrxI2iyx9XEuQSuA0KFrsyoUxScWNk6tjje4iHBCQvNoPI0SxeJnrhkoyf1ECw9
cEAEB3uAzgOkqlHaV8hskyYkPj2tdH0bFhOpRvMfR/DWashGYQh3P7M9NlV+NFBF9b0i3CiO48Oc
WzpJ7kWYypbXUvmx9GKYLvd/UzNy4gQZUjPZhFLrFwwDat40eQ+kdOTwCaPy3olkJifEdfiXA+bN
MB7sr6PulsnKFuCqvcAmxvpyNUJTY3T0xBNCuFpmgPJ+u3cr5tC02P6Q4XTfYgnrfpigzN0wiZqc
9zpn4Z5OXbrOJi2d/BZ6YF4ClDnj6H4KBOFkCu37dMz1j9PCd8OV6Ab7jdprGHAYr3Gp51dI3AwW
ZSJwmt9lAfT2ZaR6TVu4ZZxficO0DFLl9inJnKffnstMh06q6d6aaY8eWDTVedatZaiJTYg25Pfh
Jf6fpSodlOE4WdLnMfBT9AkyUU8eHrOfOIPpLh2qm46mt48LSyCO2vzaV/+1foqfECAeYRgWzC1K
SYyYw6g+iW0lGQ906jSeFDluV4rUVMqbJ6ODt+7mg1ft7acJVT+Ha3rdsglwY3wzeaqsryN8Y8ja
nMIfeW+qWHrgmLxRN5yrhaSmkTHcN0BBV1/1RqGZJzhfgawTc6khURazbtlir42X5bN6JP8Ra9sY
aAtzjk3x2a1gVfaF/V4oovGBSa3qWKL9kR8sYzAR3BA7T6jENdWYEcm3kIiTpe4HVY62+eMJvR/2
xSUh4mnDmrkhODHq4sON6xh+dvGrsQHMeRSCLl54uMysn5TdSpbFlpo71va2NHWbuUfa74J7UIVc
JYywT7J/g+R4eWsoBG1hnwLnjHGxuK3s+l45JwZtstWsygOJ2L0cLByiWK3mgIy/K/d5sbE2FC/W
/yUfCfaIxOWuQd6DlRPNYcsdO5rAf4Wi2BGfuiQJhOPhl3i7z/fMl6LSdCM5+9Ztk2J4C4O5USsX
duDz/HV6ybJF3VIcUwxvzZN1GW4txU9qS/H/xgeyUDyJxz7itlQUaQvuprhdVrIEwD8Gz3GddpOS
970/KkQe3V/l3C76jBLLfY6H2etCkkiewgll15ufFFGHBHjMmJm2lO35weLwSpcWvVUUezyzfsot
FoTTRsYNXoLEo6VVjQh+Ltfvxgd6tDgGruyUxqCwnsr5bYlPoAj0Pmg2WwE9p8Ang7dIRjjCAoiS
XK2NPSs6wd870P5xkSMRM55T6oPW1K53Glb85py5d4LkkEK+6ncMlCroJCCLDpjP0JqpMvNKGBI/
4QZtG2HmSY9iG4rD7Pfu626Ngeh7SY2Dcccp9ryFuKR6qrp74JcHp3sJqDOiaMKZf+jwpx4v/OQh
ScMHWK+0MSIFWdz9smOGh8QdCtLRZxABQrh4lGya/KKuXVNqWlaVvvwOa7OLMH75Wf132mCzms2F
VebjcmNnHAMpny8BFKd++tIlhGf0RprBTybGjzQFs7FNlMS4y3e+YPsKYKmXYqrBVMRC7Qe2Ehyj
ss4hYiI7uxATc7q+gvr7ruLh6u0T9AXXz1wwqoh2c1UXS4zpwLkDfLiQjKZEFzN+kGEoezQ3NHdk
L4+3k0oMF3KVcrLnSQA5gsiZYLa8boNCHv3yBeckAhViFwdoWORRfYJs52wWdc2hWeyfj1I3Ksrt
qkD4Qdx41K47D5rPNTRz1DtACJS0671ai44gQJSqSKhpEtAyuVyvMfycmLP6KBVmZ8wox6Xh2pS9
4LAAzpItfIfMycBPKAdcG1e/1stCjjIiY2u8FyHRNrHOomO/hxBMmSFCd+8l7OPN4cPWnfKAoPvK
s3c5H5EHJU+sFIrPupcmOirkB1mQ11ipjJavc5Ophwn86zq4NNR12SBkipgDha5QLp96DquyhOmY
1NNm0F9HfToBPm7M+XEQ0M54z9w8OIUsJGcNR+k1bhnmKAuRZ4WrMTBWEUu2H4WSXhTd+v15A8it
DwE81YHeamfQg/KDykPAJ8058JNSIi2ERljjKN8GIrNkcVlKHM6lgiHIyWKaRNvulHlaOWHRFeEJ
FyX0Slo8GuYSf5IEuKu5LWRhTRkn1q9IaUgxjWGAlxRzE5rEk89woewIx7gItawC+r4Dh8YSyNDD
6u8hO7VdWWkGNP1cHYhuaxNGjDkCDRTjphuAg81c1zGrdiVpXIljkPxZjViI036Icr3c3h5Cxn05
EaHFtYGcdgk+iYpYF4mcvjUeBx0L1DuqCDrhtKgGB67QiYwE9kqlusoQDrTE7GLebFoQXPE1ylh/
XGB6LyzLzV7BdwN0GaWsYZWppMZlpzt/xm6mBzdbc79TM5Jya+d5vk4DaRHCPzujVw73+HMT/F6v
8LS2cchhbh4+Z2/BRtVyBlT9eam5q0JprkPQp8AQowvdL6LqBGnWjqdMm3Sx1P2/+o21E5wxsB+v
pEq9zacdGnmS23+SQ95xhetikaAUn6U1zzDwObmwyUIhbI3gPPUYc+3I7mHL300ElWj4fWhiN/Rp
NIwlih1VNf791MDvHd0D5cJQ0V9yHk1w0MbgF2juNaPsfQaLYqcf6bXqwdPZCsNWQFWgfm3XTGVt
eBh6eKCUMMasTNwB24m0CgKGoQjl4n4jNT6SpycWTLxyaJFgN1vA+xnE8DtZQCmmLK/MwcQ+APlR
tUP1OGYCCCMKamZYwAOlMBekG+mep1qc6es7YfB+z4XnmG20LUZlS64E5TOJ2HGcdSacop8uthZB
aoTEkXPPyrDwmz4g4PqCbzCRP/05TmOoCPIL2fqImlkwEL9MIEjZUHVTeZShs/6i/KJNcCeYGP+u
ZQmGXismPa/QsWZmEI63v8l1QLdle59V2Wpjbf5JifUZyJK8n4RNwQcyEJDfypzxikzbRuIkgYzP
mKfd+fFrZ8PjMWZE+1q/+KrKpG3GgisnWKL9bNIrjpiFPqXPC6FY8orCRZ36Ve4YBCyedFH0LOAK
VeZDEc+CHH2L0YoB/3pPeR54SQxXULvzV7ubCQoOBm9OqJrF9r7IYE2zNo9rIU+r+i94jayAMvrb
t5DR1cSK3yffgktOHS/2ky3OJaOBrncmA1fxtaVYlnUrsztZrzibo8znW8w7rr2Pp/GyNXtOP9II
khQhVWcRkpfvG2CJ13ldBjFNxYQg6UTvVeCoQf0TbLrDNrKnNxBZcKagZB5H1itApNLmJbYqXueL
wSHIac0QFP1F1qPcddszsfd0gAf3clj1R2OWYat0dQSo0k7h3wfSawNvrO0o8BUP2WFKDXl4M6Xe
1N4wZR4noYMsrF/52g/ko8DplTQh5XHVX6Kq0smWDvEZan58AT7ITXr3l1wwTkEoh/gWjB/EfNQv
4plZXGqi7lDAiWdBh2lU4VY7duTW1F/I4Lk6rZD95Qlssyffh91OmjHzPJoaavtkacz+G+xfHPOl
Tc4De4yqa9BXzSK3HuTi9wDGU6yf0FwlWPaXopD7VVD4z/ypxj1ML/WhHemudkGQCvuTidnrY7+p
riBpqyGTc377Di/cJKIZK/TAiqMRwuUluyoscGr/ysHvVNvkKDyKWVGctwqsLsc2Wm486XHrQeDD
yjv6CQz5iVlCSigViLH2cUJjCVK/73MURr8ZChuFw4NfCsKFfhHm/zR/llyR4YHewzRHLZLSUmZA
AXL66kcyhe46XvNBhrZEbRVyJvLGb7VG+iHCezHpZxzIwvJtFSHO6uAM/P5+1R56yUthSsE1u++z
Km1h2fF9lm+2/hg0mv8BI2TAxWMBHYl2KXSmc4cXclfubxEaAzmF7AmDzbsLHGf1lKmPf0/gUga7
+lC2JpvKj/YZQ/CfKl8W3WL3mnJ7Vmk6Dfq7trLKZzygTawMaO2LMy2OnNpqW4EWyast6pG3clq8
W3wkqq7vEXuqfcmCHaYiCaAGuXx5SnISlvbmScF6n4Av0Tl/+q85xqCKf89icYl8egzeaUOpL41m
EUHezvPTev7ngVbTLSBmo/bHlZXb1d1vNaDjTonqe096844XBC3xxd9r7zPOqNYXczxvwj8mXi/W
BsQTHY3ZALEyYwm2iMjd5E+DkPV4zCam6R+0SaoOAgFp6cMNteYxe/xaxA2PqSQfDHOA7lZKgKvX
+6wmXPV7C5bFPwAEauvlQL/bd3lJNVlTSjuVuqeZ9Z13arB4LNPWZzu7eAnaeLK5QaVktCmLL2Du
p++E5tqUFGHkI+RXwfBInJHuoKIwFxRpcHHxkXlbxF4/zo3IHfHyRkZewpWf6U0j6MS4NIUJXbyW
aeaWGIDfGxIreqON3+bOvQDLoLoKto9kJED0o7hyaxyx8P3AI1tUhVjzGrCTJhsrmyQG4glYzdBa
++4hLYerpdtLO9+oBayp77fDQBV5W71TzeZJEEp7ESySZPV9rK57ODM/4d3Pf7ouqVQ8lApb8PU6
ACaUFdgEJaso6IB3YsGuO10FtBdwWoK0KoG+fk18j5SLJm8JEV2ivZBE0BFuTQU8+T+v9i9ELOI3
wlqehZdrZUqYt/cc1sSF3/T9DFpSkLUlpRjaaUyZsydNkWea3sGvkv1QLXp5JkIdcaFNPPM+AxuT
CBNheDoikGeZKgKyjI69UJr74/MrlDelvTYhlWdBdTHVa6G3DYgeBcTaqoib7JtzbKqYnisPufv/
J3fyPSQJvkZUfuW0956jWtMz3ve7j8eVYJ9QAHFbM4ljue0ZE4VOSDshqCSETWi6w4xO8EgXM/uO
rjK9MvOFATUiXj4AZY4UVPsy72I06/el2OGwLwEabOu0cP8vrrq7yhtK4p+PMkIuTZehn4Tu1tlY
GU5FQMeQNrhpZUZSZB7MmdA5X3rC+Cq5h+Qv0LURLV6weivONkxtou2V409x6V+B2C+8W3Vfc0L+
vK4XGAdUoiNCGXzjPxzpdG3s7hDGNK+eOXk5Jun5UnZ0Apuh5VRY8+212t9QRCk7gngwAVobaN0w
EPHnEUdnN6RITHMIYqiwG95H8ZpL+T7hfpm4LLl9e79Q1rHUjmCwTnLry4WTyOM1DT3KAUtEPSIF
Pzuz2L1l2sm1I+qFK4UbXUosD36Dm3WrR+4Ky8xTAVcOSKarsbw+zksGQZRtTN31NF+7foPlhnmh
/kuumfRNcgEdjvJQNxKFtpNJLDOxnNdsHaSA8VJXbMk5uC+AvgXNn+i0pSTKU0jKi+NgJc5kj26n
eRk+4w/ay9EYuPw4ab1ZW+RHi8btYFfhItsPkbET9E3z/6mloLiXzX7Hd8uXgxxSq3tl4+VGGEb5
sgdzkS/h69Yj6ve1DKPQW2CVLGZQQ7w9kewp4I3XhM/Y1xGyJ56sUIEpMQCtibup66cHkIX1PX7E
uGVFZBjJdWk0OVDdaOCrnYYZyWMsA3Y+0bebleS1ZBWhv+VmpYFIHwVJDi7DvJypzEzP1jrK9x+y
FEs7ujFepELuX38jRTqeO9Sc2c978RvaHtZF7U7gWd8fshv29M5SJQS4fbQ/5/nwVy+Tdrrx51Q4
tbeE3+do1MLhArPrZmjv5hkYgs8X1RqHQGdnnwNhKGAp3RQRMJoJ0r0SmJ5mLaLdUCxhSERmL9U1
FXnundYqHdd9VIEqgTUhbp4vws8bLEX0gMwPB1x+ULhcfl7wsbglDOUCen0gsZM7iI09WaF23FUK
lneEaFEvtHP3bbxxmJMUyRH/NWA/x/jDeCAImtJ+jxIqLgl0O6TVu5VyoYNXugFVrDLGNHbL2rsy
nMHlIYTiqTFeGQsBvcl+kaG4H6MHfOnE4/CpC56eI69gR8HiNe6TqSxbQKlgCp7KmxfuOIfdJf9C
B8Puxg1fvWqbLICeCkxGJ2bHGbk51gV0eCKtwlosZTWooa0CGiRXDbxK72UI3rqyMLmSWpUMIDfM
0n5gxYgrXbXECJUiAAFgYL4m1AhmDG/OqEkIdcfDcASI6VvvrVvFzX/HSgArKEs3RFmMTTj8l2Jw
60uq9oBUdfRpZhEj7c8k2d01S9LrZrsmmx41RPp36kaFSrhUvwAdI/SmxuqaIf6tgSj5UvkPFHbT
NO/p+yCD4unduD5w7R6rCQ50+tLUh8KBlMXTHoF7harLw+oMjbnE2NWadSUSLuAludvYVY9cdmQ3
9f4C4zYWMap4rmXT7z4S0cQrmy5RHhi6Bd18yjL0/QkpyKQ6cTyPL94NC0OU5ffpvo49ESaIRwGm
ofl2wypVC0nNsZ4a30V9dg507Z+P/dECjOWmn7yrDRs0Bxh5jm/gwArL9wgaH561txWvMPS+JxWn
CvKHAd0X9upZMcHzftNsjRVD80Wb6XIGn8czcgDUFfQ7GR5zmykrkbm0iR6PEGDtonYyQMkUBeTw
RiYNwo+3h8w4AL+PNTyde9k5G3UOXvnNIys31xSFw3hLJcTAhkVbsHiYRmKDv7oiW1si6W6dcxQP
Tt0z0zBMIn4BdRfMm6sMSKkSMvsho6BnxuRSDS66+4+YVVgv9DA9YBxqhysyHvTCy7/gtT8ebNTQ
Mi8wO36WI4ngZ+/nswB0BVMENXOHdfqAQdi0oZaOe4QFeZ8FNa2Y4H7/KdEsKvLQ3MpjplSueOBD
uCpkfl9fQEWkidGWSvEaeXp8FeDDirTRyTKjyBANj/3b9VcOI+w10l/hCkEAFaKxYSbzeTvRVZgh
6SfLSVoSl8TVmof9jj60e+TChnzzqYNkytsfF0KWJ29ntP4MEbRqisWaHaLQWp9mBusnRY9glD+s
KvsG3WH2inv4tmJbkXqXZmeHEIVFzQG8/Z2pL4suPo+/PEE8IDp3EnPUy/EumsYEVTAtfTCxt84B
7I1rrEsxn1jvcjVBNd6zUEJeQDuGx2LiJBsa0EAXikidlvFMhmQg9gT7ykuMJxzk1472quL7pdFW
wEudMeJIYQcOa4Fn/9V0Iq3dKMidEGXiEKS+MjM9yL46tuR5gtUh8vQ24PLX7r6I6dblGPkJIKBr
XawEpRiEqOHAfqRkWkAFoZBjl7M1ZIMv3LSPHcGJ0e+5bwYUppaM5DUo27ez9Kj0EL8aKOARuHxA
ZVhzw+7C8f2lmEF1WsLkBtUbcWf71arV/uegWqrzeehMeK6xJnWrlgv0tmvujqeBHxDtz0wc2ogf
0vrQ6FXFysIbS9L6jMsK/4RFpjYFTDRc6Qzzxb7gpAuOX2aEbzAeD7KpTngVlcerkxR2B8VoKZZ6
e/di6lYa7NQRgsspYOaSOgz+8HrYl75yTGqE00Qna1qjuxDLjSw1A4geGtsDlr3yGVr75kdUCOrX
Ye+5ujaL+0iuzr8CFYtDIgRjjNyTyIp6s0IO5cHx9/IYCg26YjNmVUMrj763gRbrwXwlc2/JjZAQ
2QG42BJWVL1nWKkoccGdba80yaQCyX7/b87i0Hhsx22hMocQ0JJjXxLiSQzI2k46/j07z2XSHUtC
xvyQMVX/niggrAbrFiEnzxbTqV+gSNqI3X1olxiJ4m/fuNv0Ih9ecXrbdkSSmJY2lyDjovAXUw/E
ATzmraUDJS0AsLmYWI6FMCboLW0e8OOAkayIVZnuF/0CDN/JiIvAIKC38Uh5IgPfe3a1FessqNIV
f8YAT/nOfxnLdrEA2hIqODM8+lLsQbSB7Hgr9L4INItZxUL4yyHKUgWk2Oc33cDeD6UvbmrSP3It
ldC/RfWkXXKsJSFyNVs+a10dlHl0Ay1yTOXop1v+U4m11QM+hlEDUrAb6D8uw7HOqDurHfthM9y1
sSU8onDc2Xam4pWtTxi6rQ7HhnrqHoyD86g64mU82rJYzTaMGovA2yXOdkr9VeEoR9v1v5JgnXkL
LSU53IdSYw4XiB8uegaIm5vsxTGGeWS04YMT0qbY/fG2aU2GkMqgiFXOXqCsPG2KI5lULgN3DL2d
9S2fAAnBRavH50pJjqycMHKowCzMJ3b0asKYA4crYV7WAFWktw2aonnS0spM4ilo2IzGFhifHN9/
yAlGnotKFUU00VGFFVw20eGVYuj4NdbTv+Dr1xdKMLov7FAdcSOoUae5yxW977cS0GFZSMIQAJ+h
85YDycOksVD3u8xE7Q8hOOQR9sZPJp+5YUbgAYepH8YPV9Wv6FVArcOnzgMt48Lx/e6cPxF/lOIf
I3r5FKbYqPiXfxjWOzo45NAH0HEV34NPM5T6fYezY7M1Ea3cI4Qf1XDpRw00lBKkdJb+CBKHJAqC
g6qxBTp0jL64FDlH6Fn4/oCkaKIsZ5STtw+6OY/Rx3Y8jI/H9Y3YW5ZzPWsyg5Q0WJzlakiPLwk9
TqEriJwDcYgTT5ieOpf7nohN3NTs4H/QxSybZTjSM7yyhePcWGMuOmwL4O3g2sXrw+AfZ88pD4cF
3d1GAFcOfzG097ZBILR3u744gvn/Olclf1qYFpqJ/R7pHQI2vjcR9asvbKvCoqrYu3FFkD4NMXL4
058GqIUmpKah92SvfSy1iBaVV6r6LnWn5j/SOspErdy6hAcIUz46mptYBzq3vSUemxJq+JPQAepD
AdkLH5ZwKbRSgitj74PdO8DyTsREr1Ym087QkYsSHgUG2YbyHxItBxChTEdo8IRNFXAwPimQtNvu
oQ9caKJPeSqOs/bVMZU9QFR6lO4bvIZfeqkD45dy/+KsvD1V/Bm9F1EAMtm8Ux7G+N+grBOL7vFl
Kipl2dxv4KJAixg8y3ZHv3NXoVbIuCWExsqzlNuYkP4/DVLthzA7gpSWGGescMCvvtbBbxDAH2tV
AjnTx/ltjenmVwYvS3k0WD7VvQcaR5UNOu5MFRR0BaOwDdXSFYEDTOSX07eKSVCkEbzuh0aTl6Up
hxTtQGnOhr48GGtb2WpcLaaeUUBwZFGloEzVzaPDR3kTPbyr8DCg9WnynXhrmt68cjv765j7suMW
WWPCLNMb6KLlpsAQ+Cu4ar8jpjECpseN7TbPd5y+Hc7ri0UsWVcn5zDbxm5hV/Iz9a4Rlbftqged
NXx8JzFRtCFLCBDG4ybeJ8xCyVrQM8mspr94YQ3yPR/fIpJdWpFpzu9HOc53tHHcBe4KgbpucUg4
0+CGJWVeX55DWyKQ4TsKqkwSpfthT6Zk8tYYGxnH52rychFcBxqSVJomPUeXMFuqqIH7Y/CCLoiI
7AeX+FW4uj9aPdwG6POokS59S+BYKeAsLSfUolHg74DUKqoUx1If9sGty1Nic+iHqTHnE/2EH0JN
NwfL/Lq4WdrMqlOY1fWdMq/JZepROqqONYD6YtUdtD9vj2pVDEt8Gx5fxC0Y91b2DpUlmE93Hy40
PmhKnYfv9j3FsxqbTtB3qHMuJoEygXx87EURFOZ4/7lHeyQbuseoO382c+98PaahgORA4SLd92h3
l5CLOJ7vJ+1cr+Qv4f3O3oGhj6LyafDv7fVGuwvDsYTrl0FMVTBMKSNTDjCU9E4FvqjdoOdc4/HF
7NgEW6GbwU6vG7XMdVZTio+6Sm0XMYnTqIvzdhXb3i0914s/wNMhCXnn05hj0t25ljyom5nSvCsv
1xWzHkI7zN65zKig2Tpyw1jYLTAbYQmxMZ5d+kQtvD3aGRPanB4+Rab1q7cvV6Aahalmz15Q2aLg
6sr7jfDc+NASDVnPlq7VRVUinmIYcGB7TpXlVOb7mDmKaZuE5bK1sSSzpn7263315JywSJ3v7vNx
KKsVHNp57u1mJNAxWiGqtB0oUfmQXNL11lHUiSrT9OXF+R2ujLkGUVjh8vcxYWcM2PtlnvuoLHQf
wSe686RLP/X6cvlQYN4CjeH159RLPyo+0vj2q6hB2wozjiZyvKYfu6Z9anPn+PAnzswJfDW0FxEs
ngsSyCmh2hSrD386AP/9ItjdbuLusRPkgZOZ7LP3ga+QRMpSMOncqD3qNkCdt45EI7uAMW9u94jf
A8qygu2i2hfpNQYrxSyXyyExfYgxWHODnsDRbCLmcCtW2Gi8bVq36rKInEydjM6mfbPo0WjQ9kiS
QSCMSECyJuKm3P+1hYFOfOmaU7wDV9O56J1nj15TuqYpJg7mRG0FRG1eSBG9J5ggLGwsv/2wJhqv
4RisoaN7iV3zAupm54mglaQBGiB3R34ngjjWb+gKYQpnT7INaL2EmeIE0OV75qCffFnS3Xxp2v8s
dqucgHhLEL3XO53KGuxZ3dLXJstnydnZkcejSX6jhDiySnj+/4W7jA40AZYTf/Hdkl8lGL+d10Oq
J036bN9x9W+r0yGBuVK2wsdTfOP56okuYVn5yDL+w70HXayokDGMIkZs79vRJAk/3YVtbwVmkSpC
+JMgX0o9QeXeKhlIP0OTUz3HrNdcyBZEvLum9hmM/tUExwM3fPQKgAbYlIYgl0Qxc9d9fGIMs7Ja
LxnnzDQoibWpVx7EoHsUahwS0tz7ZUtOBZ16UGe4GmO+qmmyZFxyCip75W9g0OrNhD5bg0Tm6G8x
/RtBW8jTEhKklKI7fHjDrKed9LIbrqvJSI3zNieJ/x+GFP1s1D0D+fZJDtoV5mLW14CnycejknEV
esN4VRmUSxRc1w4I08W0yl4jEvWKIPO0uVervAC4n+VVAGbdCOt/8uuirWg4paHbejUbXDd2lUit
hdVh2y8FdwMu4QF2SO+TbacyGwo5TgwMiuo4IK6OHOvGIh1DTOpQ5ODqTmeuTrRzk1JplnpdzdoK
a7dYclv+irQEZh+GumDCDS5fjC7S50kWZBPXSnmXo+lylatHli72+k3TiY6Pv9f/Gewp6f8eeN/S
mBujovIT2UV50E3xGIdpUNvAKOgb6bf5VpGHJlG6TtPvHcMM/DniRZ8BpETFtloGBJc6CEYD/wbK
MIsDn/K747lW11MQ2NhqnCET2AKP1i4q/oPG0zQsu73p/71RNnvZJZnt5rcA9v3ixz7knlD1r3L2
uMl1nKO4QyCN4SZSj9b4OXta2pDjy1fGoSXA0UVrYCSAO3j0Bxz+MSMsfSp3h30TypWrGcoqaP5v
Xsk5+yzYe3JqAnc89vimVmpteAG6Zno+pLHv7BmoNBye+lumzWAJsPgF21dIDxn6NvfCjtLMvjJW
CIBqMw7zskA6SUho9hh/46Az5wkG++gTJVwNaqnEfYUDhnwme4fhsUsedRXg52Y+Es/Afi4Q3h5Q
jtStuqD0rdrE5zTZrYkEjr/11iJ/QlNM5Gm/BcUbJtIUPaR3ENRkxBIr7nqA5oyizDJuHrgPdXfX
/ANjxZdB7MYBo0FreDTSWyQwhSiq2irH151a9+2w93cPqv6Z6j7xVwPMJkn2ZejnvwfUXH4npbZu
GkbPY5wrbz2Ll7qgSJdWGUUTBg/GLMHHO8fHct+She0FdUlmB7mBYlzoRsofAvORh9iJF2kMql3I
ycPMYkz+PNWwf/E7j2zbdATxBU9las6CPlmkWrfNFWNtaVO/C8bYR9ur5zjg8l5C99vmrcOD3r71
3/D26N4PIssx4RcvrVPvNYIRjeWCd7CngjOrzyns8pJEcoHahGeqslc5OgDJbSFZgzPDoaKUy8Wl
772RC95Q/l7Gr2v+6P+CWHxBZhph3wfiOURgbYw7jlkcQrMmhYSza9ysMpR+xdRJwnALZc0phAZ9
Wo+Py0LiLQdze8fgFufPLd6xaIKgKY1GwYx9AFppAPzFsnRYZjTU2RB0fPDZU2k9Vm1WKZUdxdEi
q7ZU3M1afdB8m3sWWUSHClwAmKhEyhh8P5t4YBZZEFdknVJybnC36Um7bVYzVJ1TyRXm1RBsZSMP
xxPk7y3dsHa7WYVvzfy7D2mv7isKpxiy69vFoE3wt3tEKBhTu0KD6oIbFcBtlFZIz/9V3GkYGc8P
3WMEMFkltHqF8WSi844nzqUDLXdzUEdey50TP1XkPuP7WhvJSpZJR7P5tx6YSBT7FHic1t27oOCe
slKrL29O8OrCHYX4Q6G6O4F8k0Html/ngNCxbhfyiGgAzs4gMFNdJ9W+zmw+xN3TbUvS+IHdJz4Y
Wy0k2gGHpUEEz6HOtJ+0jJFm8PMevKHV/K026jRYQS2UrHPeytRuDDiww8p+Pn3a8pFZVOgrtr+S
bnZc1vsl+ZYAW8aRnNm6PNvW/4hwjVnGZVaVWJvDJ9hbd0YV8E+dyCPtFWyuA1Fx851jOgwyde39
dkhLxe553Qls9jkvgqgNhvVWbZ8+0Gq/Vx5XDfpethYuLMw3hk201wynbb7w3ep6LU8hndRF0Ybw
ucWiQ2aVJHWs6p1WhQhTCL8ZmT9eedb3w+y8iQwvbkjU0Nq/H00tEkUb22LvZbSEjjySSODhQXpz
j+D3HRe2K7Gmf5MBlsSZGf9q8KH7KNsm28ImJvfqLdiKJzSC8jbuI0zLmIi6fxn7kLpoLQE8WbH0
8mkBRu+JXR8I9I0kRKk/fYCmH+ALjq8Rva+PoyknPUqi3KjLkrE2Xy7YSZY8usz1LuSp83dZ+b6v
J6zCkyN9rHmFhl4ePEtMpN09vy/MW4PD8g7RHaD6J80ETGxzLsn8zz5VD+06OCPlFEkSUOrPzRnw
OTEcUdf4XchhOfHzXBOxsAgIXGbtfbVrDZvSOAankRQ31Ea8HEfJD5/y0guu4kZUfkVyU46MQ/y3
P1wC3VOFUErqj+eKatM+9/8DB63xoRzA2yFaIngBA/DTWJmTt2miich0h1wrGqcwRggm5KWnETHQ
kmnozOKOWF3HVKuONI9weBEa1j5PkW+px3qDVl0VrNtZK/z26sSDF6P6I4KliBhHQgjLp9wF4vFK
nWMbVx1wKmSQmDtnLG575qkiN60cTcyShdvBXHijrwM/UeCARdbc7N5NqwJTQzBkZ5jRHYPmvxjJ
pMwScuxTrYN2rZPM5ywKEj/iSZwZmv2k7/D84Afal6qJxAPDxzfjDsbz0VUF6xCtSzs/yH5GThL0
p0PHyu+A7q14Pypgoi6pRy8duJ2aLF+a4O74vvvALsnLkJNckY1XyXREBxR/fIc+gmXzXDONiU/V
Zjbo+iFMM+zhkqJVWehEV+IlfuGoVy5wAQ5pw+mYsBCBaQmaIvgUbwXEGWKZ1E1tgJT1ScLcgE8W
SH3Xe/NnyQlr+rEF1/PE2KpCcc3zeBw08jJrswaC1hSTWRQiYVaHPVT8T2atONVrD9TILqO8qL9R
MXoXgNQzVMa2GOYShq7LGB5ZjELKlkU95+TqVn2G/+iIIu3xtrrUGv97HJQuEtjfIKaLnqViXMY1
EBw/+F9xVmZZmcZH+Hu3iQwnSRQXfexac6ep/NWyX5T2K1EuNVJNDI2vhB+mCtl9byggCB2szM7w
o76/owwMgg4Khk7o/nyW8uwc18C0Zg6h4ed49HoFg4blB/E/IXcF7UnA/yJMxWPzRX5OPpSbmDcF
2m22b40r+GKYVks8cQe9L3N8BxqDg423XJ3DUhjI3nI+z5Ls5K8Rt+8/eg2vj3t1fYE/JZ1uGGzk
LdCYXuXmkNsf/OBBa0YSVb7g0I2zf4/5fBtDrMpWADQjoYyIr6JFK3SSWcSpUWcAqc57DVbXuvNp
HEUvoWPZ01Wz0vR7sFVOpifZtiOJxF1qaMQzBBndflSQldVFfMFxriq4m39mpMJfX3vwIgzf4M1R
ZbP51HzUWkw9yKJTlNf8R5XMAVne303WiC9lUB6HFTAa6mJ1L0x8z5RuVqykRiKgvm6EzftQP3aA
GUeI12ucOHIcN1i6/PFEcHG1GncMYohJu2qiSPoX+eRbIMblSdYu6yiZ+SMXoahb4IZ6hpDEcTCb
axjX69TMb4HTLwxRBD4w/cevaVmxf2xEwmFqFwe1mSonM8eDZ7ilydke8yifJ/u3I+bL5nhZbuMH
sbbTYCzOawyQuXkPiWRan60Cgv+k1tegpKiGkGeuT0LbfIkpH58rQA+zxxgtYoNb2gp1uW98sTQf
UNYcbP1m8YPMIrjRgc70yn7t1UPmHyz82y8bzc3kpoVlnFpEpWURrO+bC9KXzlY2cRgKk7XGc0Bd
Ud2CkjoPEcRMC0tWFRtEEhPMngUUCc84+ThQlJv7gkHIzPRzuK0uo2LPE3/PITX2dq2pnTx78tH9
055pbuXeVlMMfWQecgeD+teH1Jl5yC3W08i2DKZwmdMSbIj5IaQfF+O8si4/mXoX4N9m0di3Y+XE
ohG2gfQzFzW+YFEYAr5FqMmk/EBa0qBYXiA7nP+D9KLl0xEtIpVzZcRR2FDOSRa0IW3QODs8eeZO
Rff0dj9/LPONPHiMC8t8XlJzZ7bY1Y3bSK6Eb1bJwGpnSr2kdvmTv6uuL2zwMFgO8F3An5x7KFvc
APvVUTxoGrXNcvPnidsT0qFfxhxB+mM547iDB+Qq7ut9q5rZPjcNe8gOy0bA7pIBAQeaPvZ/0ndA
LRZiY1c2f2+jiIkdAH2KtKAx9P8+9ckK9Ac5sq8yFdW5bmdj6pAF539i8bugXhHeifqx3JrB9o+3
ypIz1KBkJAOd+g8vyX4Ee/5XQnkcJDQKkh2671Ol3QQUe3GW2M484zs7OsqszHxlrnH6u/4fa++Y
FUcxHL4PlTAq3LzZxiaglV8uOQ3pRJ1Ce0JyISe+Vq6tXLVzuFc4GOiAS9/LlNneQv7jRbVkMm85
xtRKXpYAREiuqZrsoUiS90q+0cu5fNtEPTuP39ICqUMJh4TBD0xHOT7IOcBvTLd8o1qplF7fDoJc
YzBg6R+qTB9n5i0VON9qv6On1YVtAkHrsGzTyPNYZ72FL9wgzNltJC5lJ3yQATKnVDdIE7TEbo/1
z0IUOcL3DF3sY0V/laES19BD7Q5s9K3XYVTVrNrXra3gFhX/PFPXvS+C5vgyCzmw1XMoWN8YGyH1
wHG3N88EhpB+2FLmSQ6EsWT+R+u+3z/yPGTFU00Sj7Ui7iGxFa5DCISvbr9rg//4bEXbZFSkw/Zn
TkA9lv16SAf2zIWbJWgxk/UN19q4cCUHSGGGssF+Ye6eR9Oz4ZWWzks92fLfAMpy4at8PEYq8T/t
AcyZsefUJuyn70PJbcZftFm57X8IDelAMTtH5H+sRVN/Xnt4ioIeFmxWIeeIv7OVHnq83xtKNfT0
VEW3av8nRI0UFF97DrFi3phm6iT4uXCC61XHJsTQ3YA+jZU1qmS8Hwb4WaLh5EdDAhQ+u0D+w/q5
JvGWDoComOOInUcUciwIqVsiXMqA7d+z2yfJxCDgOmB/nC1s0d/LrkfF/PrsRAlYLxk7KgUQN7Ek
mHuDlYX8H2D8Wzk/azzmj9SjMXlD56tA+3WVBlP/VjQecL3xPYUNBT0mp24wSuQcB8wG+h4pIxg1
Vh0r2wL7KTm5mV4TqnhUQ92VDaui941Ups/wu+vIaZVvPt47/zgxxTwvixUl7+OGh7s1hkbK8A3m
ncFrtA/Da3KxNb4e8KGALFDPvOHW50RX8Wq8OFnDWLLRtWoshH+DpxTDCb9Ypfdpy3qoZw2FPXkG
y5WFx0GuxZK9YLJHJlfobEWSDfUDu3PXFOJSvWCECAHLQjBqIEMtZT7pDkAM0cWmAytH7mCK7f18
SYplf1PBe8jipi31CvQULWG8MyBPHInI2Sf9IcOFgUUMUNYeZsDlqHIaznfDTzI9EGjyEQLBgOQc
uwdseOPBf+TpswqGW6TupBrkSy7CRfqfPn+jsz9cXxs0gTq0wjM6cTnsej/NRAFTQ/day3WEh44m
SE3m15OS16B0isJ/xsJCdMwHa2+drDCwRMfEomAJdWW+ZhWsZ/s5YgKGJt81L7Wc32877JqbSKH3
udv7eEJ3Ur5trM2juYvXiDXC7PKwdGjKvqSK2+Bum1D9gxVE2FPwT1akiHznN7RCVFvMHszZwMso
CglsRGQwk4EFIzyNX2NJi989H6YaEQgWS8bAns+ZEHhUpwuMgmpg6g3LMe83APWX66IkWSFnu2Hj
XkX4ClLT9yResfbtNQO8MPaashZqvW7ECyo7w/Kb6R9W0zHoMaib9V6jwsLZiIX1cyq4xztuYwit
+gk/xVTLfKGC/Qre2yxLRI3sAR0PrIk8DaNbpZNt1BuPSsL1OHlf4o/e4NWJadROnIepA0BEhd6q
VX1j1+OB/wY0t97kVlA47p1Na6FvUkY1UJI5elpQtAyKgBcbKLVDWO0hxXBRWQFxFMfMa4yo1NTZ
kvdf1HGNl38IV8TaU6Pi2+Ap12bDaG5Ey+Pz9lImsAGv1B4s81g8j1gD9HdMEzncJzacQOhu6n0W
cSe65oz78aX7ytNmxr6wj65JpvxUT7mfECWzhyeyPpNNIBElG+iB1UShoG8IjSkxZYDPEdPQ16ev
O4TmfpGfv/KVyW6jhJ7bThiwrR9eIY3zB4J5RYj6GA3cYk0TkCMP465qad+e8R+1tZBrquDkdNQK
GvQ03kx+G1Sc75CzEdhFnt9KR1OlzrDxK1QKXQzig75Rbmw9f0rhpzVXy73ohZvLHFS/d6ljGbmU
C/T7No8OigwfVTm+0iQ4xCPpaqCdR2wFzRI+gTz6dz0MEJpQK9iCXMwclBnYLGT1b1bsjyaQe+Et
vKrhbtD6r3b6qLjh/fO6qcUxW/EuPyGH1FpQo18XcU8h/rIgVhN011XWdu+3xHjTXpQe8PUmIdh7
zpGEMkSvM65K1mECf3ow4Gzp3guAQHkXCnSPmf7yqu4uvO4Qv8x1lZGB0QmPfiwAcVLF0PQnr8nK
dTQcbB5yHI9jEU6A7Xf5ITInVel76ftBnqwkz6X8+FZJinY+ijR1YeI4Z/xWxSbhE3aNgDkgBq+L
OTGNaK2EQKny6xPPBYR7xKIKyMytbfv1iHWUAbxN3BtTfsFLtU68Et20o7uBFSUfaHV0TnJMXzxL
M6+I8Uus/iI8NFHpMQfjva2fv4i0qWxWjsPrSSFKgUzMPhzzi6JpWsA0GqI268todBc3YdBLIrjt
xahiH70vtTH+P6FMW9HIXFhho5pB5ilt6Fkn71ArrEhxqH1Ik/26OsfpHe+t29ciah6Y65FkV7q2
XAtpO+RICgUyjsNXw+cLmnLXlzgCh17x/mWk5UWk/FGQEF28xf2rWboZUFeZ/fSbIhTfhQkng/hh
YZrcAITVe2Se8gYY4k8mF2AroPUZcncusP8S8vxFJFKrdQMk0GXvplcNU7dmkftHLIMjSw8azhVn
PcmOi8y/QYzcO4FNwz3ifwgr3r5j+BOT3kihZGVTalrv3Riob1GNhq8PhG2Vp02SqiDJMAactT/9
24qvYTIKOfYRFrT17QUgYUfFlUIK5BE34C2sXv3VZVEARgFuVRTYQkNJclHNIFtIk5/t3UO0qCBv
IsiWLOPo//5JWBaftQklp8KX0nvu6URVMnhl9hZ9Qoa/ed5m3l3pdpM7/dgm7bcJrYv0UoEAFGg2
gRnQ/hbm4S8N4J3nBG35yT3Uubfb9IEIedxT52ypMlvHCOM1R8EUBMkSB47R5f1vJ9H77Pq67kMG
u1ixeeAleK0EdqbXctz+sXwoH+aTe22RoaQmBOxiMwiGcu0SxlFb80eyUUy3RLRhYAMXuHUdq1zz
qCWXCd1LzK0VkL6qSYwkXTGY+ZFys1c7E1xR0euyO8hQnXW7vMGnp8TRnfd34pKnWHIk2COFHXQi
WksIN1s/abpvHI1I3PfKxnz5rqzYu68mlShNzWOSJFBNEzzW+cMiXZ7yBwF0TJYIUftl5WF4bsBu
myqLXDuWeQnqCGcF4pHjP4ib6LWiB8xQgGctQdBwNs73dZ8uVPY5eLR5MF4u31Frfje5zyx3KcFz
wxS6a2cT4PSw08FqrHYeQ1yZbNb0wubqYb6IanQj/jkPR7vzAWn4+TFmlsWcca+xyDlCPdtvljvg
NvbFgHEeUEdofVar3D5dME3tdrhqYiFhDUMuDi6b5uCMU7Bv0GDhsl2yCPg9qhK7Hmm0FHSSzt5z
ACHmj94lmaw3/N0P4CItgJmOzta1BqN7hIV34aqyDodzoXOvQuqsG8+GgtC9WljDUpPxgtZpf5Wb
UszpUFe57Up8IdxZHNqbbuELvl1N2W1pBRNC6PEqqRAsOSh2XdvKjCDoaiDfhDFX8ctcQsh+xnGh
lIMgD07lScfQZOXnVhkzyOHpJjBsMKEKHSdgW47fabW26bK6uxfL2nkMJ9zZ6pKZq9FItyJAxg4M
Vpfazm0NOAbyjC+X6mAFe9sHlEHEh9Y9s6WaFnyqLdq+n3c5H8az4hSjm/YnIhAkr3R7X0nIt0zg
1E+tZdmQUIYkAD5mlTllbcRII/tkn4Nfl/VCi9LZ6qmGAysxG4d2Hyxt9i6R0Hz6bE/U+JXaxCuZ
hrEsC3k4mG0oooVIxuKOedJR49xHkoP3nRcji9O8ufmt6m4XtjbWEhEu3Nxq5rcQ1P8asAwLTFTu
YSnTg6FB/qBROxhXITXh1LANPojh3wy2pOVYAXPQ5iJaq2qrByp1lm5cRj+Gdj5Z5JgogSZ7/g6N
EwudA3S81wW59hWQfuyzi3NV1JN83w44QuAyuC+zsAANMtp6I9SHarWfWtX4qSIMeX/aLH6SLRvr
T0QTucBFqIR3SdP/uQ0S68TzHtpuxvT1o8QtBfj5HzykG/bGuA/e9uHyMjV07mJp/+0FYQmdThxa
qj/EM6CkcyBphc2l4pxAxnDcmGqHMTmFdMTKQR0XZyDYDG1yewa8dzZ0P9U+9DbKCcBsYdkD/eBb
ZUs/O7JR0yVvXfoV2VTZhsDZWCGxg/n+t6IIuy20EnhQjthQezk1+a7YIM++5+eGlVhC3tgtBRTT
/HgLsyt9rHT1OEL+Hoi53lsJr1fS96VJ9XPZwnk0fqmIMUXykdCaInbbihur0pW1FgW03Rr+8nnc
fus/BOfFFqb7BkRBPbUjk4eM/D9HnqRbggbNdbMVeZKJ9r7I9gr1SLb8L4YmveiWpFSYyCABPvfv
VNTlHw68ycc7g64dI2Bq+i3mUkad4BpzQCYgAHxHb95zCy8n7YRfyxCZq5VetUbufI1HCGcJ6phy
GdvV/fRc/vEhnf4hgvnrGSe8o9G5+icYO8qdkW+Rr1YMZfanvA7IbXbCDJ2CsDUpaKqpON5cYLhh
mLCV8o10Im44EsjnMFRt62sqiugYKu3zYv7aP/HcjeZ1khGxXWm5QadVwEgPr+QfmRzCi6SEQe5V
FPmNF+Avop/CcsmRcCQ3/c1WWkUou0yNqht1ncXc1TH4KOGlbM57JrNFBdYH1mbz4aK3oWodPcCG
zle3XGGV3RaUx3MQ/hF1DoCWOe0RVnbyXkJAaHnhZTcZ0FYQObmwUK8c8p+2R6L7O1uCwVFUlrO/
6UBPCzhkUg7AHEzZgrSyHlB+h2CKUc0mY+5hyWP2Z4ZFRUTBt4pOLczcWtpHrLKYTuALiAzGH+0W
huSqYxWKytabNxf2AlMFtUa5zy/rKr+adXJinMmOy7e7zG6oMCAd0h8ez5Q2eLKGkNySsqSXd7NK
RABv0g9eodN1XKIgnVq/gNdJ5ObtvPPOgi5RwgWa7Y/u/Dk6CtogQXdUNPa0bplgEO85N8z261Ao
HM1PG4wXr/4qLEDcd4zr2+QAntSjLfhFIsEUDnIwuZCyczDRRcFrnwFCBnNsg0HiYAz3ZjdVNdUu
AAkPKH/W/vG5icz2wktWM8gMpc1ss9/7BjroDvHrd1edNS8y792iBZ/DeGu2y71qmC5i/xWmjY5B
1xPqFF2BZSal8I4onl/R1TlE5X8XUd+Fgsd/1BUL9cP6Sq2rdeRxUYiEJ/4XQ4GKNx+YOc9brrI6
czDbODeOS5xjbq46y918bzXAQQPuMx7mn9jSnWn6EPFNXE7tMG2CmtnTUQquQ7/qtQHocTYzomIy
CPMvqN4njXKNhlCf4k0dsIXcDeHV9yEMFxtEEzbmKKUX3GBy9zZygukT+d3zREmrJIeWqM6yu50y
F6Kq0PFF44aZyh4b3DUxfjGOQVLK8G43kPRfwgjn1b7C1i/uEwkW4n3i0WFBKxyPhANg2LrMFKlY
a8gcgdKgXfns2azlXPhDutQNCPmhz+GdfEmz2anlwAV/efhXqBp1xnTzpERgLFeZI4pbIgBocg9h
ga7KCla66Xme7Za5n/mnWBo1LWqxKVQ7+j+D/vv2/W2zP2ughOOnvn8ggATSsrh9Yzwht9zHmxdG
c+QM7sXOSqnCR26DxfrInnQLiWYX3UeERNxA18HbMQqW0izADuPldBTiGi7cGEc364DrcstjIDkx
5sWHU5y6ijLVN2bsSlLfG41fFKU/0mQ3i+96Y51ltemBnz0UtO7VMPwHotIX2+RioE5KLhOqSjjQ
slmur50QhqLsRfKCQMbukRjDPLzJsaP3IO7JT+0M+sbGommEFTxvuSWn9btJnEAFmMeo5WPkWP8T
Bj5nc5m4rKOob8oEx6JYVvCm34TQ0Eu9M8+SEDH3BvXl+vlLKbS400BztXLSRgpblu+vuMqljAMA
JH4+HEmJRX8Jm/UZxMKzawGYk5Yqo4/t5pMdblE7RCok6d5OC/hWkMyeUGk5auzj1uG0qnKHrCJe
cDVzW9n3/P1fOjbnTgvkK4ZtPXOfgiW4Iyb2ZYtM8FAi+WeQsAFuX7yziUSCtUZbhZhvvorEnQKl
DCfAeBH7v/2PR4CQarkE14TMp3VpiAiq273DFhnab6ntewHOFW1nawppnnwJgeFHZ7kUZrc+SkPs
OoyWyjSZeXsgY9DbLMTfI3DrWJ/ndFF2ydSkL5ycnHPCNSsIOoutxAYmEJYVa53/4r9OfXEQZL/9
GwoP2TWO9beSmSPI1bo3Qiqgdjl+Q/oZe1GHY+hGvVFsG+1AAj0+OlWIh/oQd7TEsO4K9mc6JTZJ
22mSh3wdzqXAF6PrLZS+FlI5TQfKz5qD/W2ioEhBhQYPweExpNJ3d08WdePv29KYvRDsZoChDDTj
l0oxHHraACIu2xLBc+8ZToRHIlvJ04MxF5wNXbiKkZeYcfhBrbxXsd4I+yxMvyOb5UobbixiSfwL
7yNvgpXviq2eC4gTSy0jRZbSnVo00iZbm1LZQq0JXG8/dtlGKT57+nuSE1Y/7Azur3fnWUwt3MHp
jmhTC2SN436wu5yUTRPCo99g6ayZvLmRjuheUrifc75qfPqtpslXVlHGOHKLXpDo9WdneCNA338H
qDQ6D0tiXVCaIH3TW7+S09e8qjrX6OcsGcxMnON+MyIqlcmERn7iA42YLnVRwtxhaIwbVIvALSlu
1h0Fe3Gby6yHOTA28LZIvnTonDMf4H56pn7nHDHjqTrcmQxVLGOXIzyTYtRMY7KC8LACZpgQ6w7F
lHtcfbpwefZxbJFFMKSs1saOdpxUgTwyJMs7o2P0Jesi2P+hIkeR1jS7HjDdHyctR/x8Nkgaf7h0
cgRctmO3EcyjGO1Axj4fCtUC+jsCseay9Z5IkadE/VTI6GKwKDQRTNtYRcOU8pJ3DT//UKTDgGfD
VEylTVWsyHtaqxqAlAp7ZT+2ueWrAgdRqW4KwlQ3Eh2WX5CkqpXUyq8331GhlSAnCQ+2JStBW2L9
k4Vi4uwxkiZAA4ihUOipRQygXkQ7sZ7+2z5DMElldau6odvXGPDm/fUnbeJ+UTGaydAiVp72ogLZ
kn4UAiF8yY3ulvKRiqHDI1ApGkhn8iuaLaCyEy5mttyxHul19Zw68LUiRaQ64wuDlR5UV2urt7ic
rJnIJ6/ef4l+5kBexShw/xXRFu2oIKiEwsSfowt7j+0kuWLRCIBNhg+Q7pEcR3j8fbRzTkkOWVPh
pXQAWctCrZ91+zqf4ZOUo9Z+HjW0Ue2cTclc4vq4l/YJsNPht0PJ5B+xcsNzCgefssurNaTZPpGc
fXNsfMarWeDvt8GUUo1GGNI112XmP0+DO6cafxnXyk9FjHfzjwaWzH6SvgWYUdecpktkxWPny8ik
l9DAe+eV8D+7j+ylWVXQ/mM5LBV4H19erNyVK9TcFmQZBJ3cH0s3vsFX6+ABt+GuwSwl/OHx0N2L
YHlz5E0nHU+3wkPd2QSnxXaMUgmsEumq7UZpsVo01g4EgMPa6DsB9bPfZw3Y20x0VZL6tF95OacW
4ICHqBJKkVRwoevI0GNoG6E2yrdP9xoufgjARI8Vzz0IbNkwuYL986slKUXcXPja06Z++LLJ1qbf
rY1r+OxF+jefMnFnED8tAk1ThtNopnCn0iWJHMvhzektFX4ztOE/nr1VsOmqN1+wi+dmEskrm9jF
wjRbcQPD8++qo3KSo//AOSVk0IzbGL+e7cck85umNdXU+11QsqqxunzhynQk+yXqydP81N0BhdJN
Ns1V1X0gM3cyONvrFudEokQYoSEqlNeFAlHQ05UeG3I9QSVJNYroDtn0Wx5Qcvh+SLdpXyHNsZoT
y1q8DIKTa2Zv8XsV1OkoAOPSDk2F3iRl0uLhnPOeRcMbYCNvDFB5eRhaPRr6Y+5W8wsr0sOVz9Dh
cGLxvW3GpM8oOuD0VG2apxTDm61j0sbVAmHDLizu7py3E3rM7oLURHacjcwkIeVt6liSyUJwmLkl
HE5M/ovaUURbiVoLbwBS6PDTwTmgiz37fksvX+Wvo8srIq4yMdSli9nv4qFAni602MlSgnCRs2Zz
haSkgkAGaY1yLNgkEe9Ri9YM1qbZSDvNV+2pw66wJWh3gjzD6+ODc7zxM8zwSiBRjLg9eK1FxOXB
N83v/jACCM8YRBXFOgZbax2Ovk6b7dwomruhCw9TK/+eTd35jJnKKlTwPJLWWm9ljqs7/5xO6qTw
SzKmVv8+tKHWHASuVSfaPIPvygodBwdgjOCv8uMXecJRThwfL/p0/0GN102/ufgRQaYOKxhxmwoU
mvVaBiVITwI4n452WiSLPFOMuJzWz7SxXjMxjO94IivOWK7mqA7hMjOzJEF8gDQfx1/JjAp/uwK/
0yPOkHpSGASwx0bspoAVrdmILM/Iig7i0lEtGFMjZ7MBaAiSRhyAfwv1GnDYeQRDEl7JqJ6c6pDA
KZ3vkjWBfEDEXgxAATZiwiEUcSVxJ+CvZLO3tUFS86vfgGzxI5e5OSQWgnYM1wtTMnVfQCMhhHKo
+4I5A9iJ8LFJG061rxTgFjIM0zIyyukTOTt7nEWnYrjRRyWJGLCiP9PoLiyxK7jt1RCMU48Fkt8X
/o1Xyd7HpBIVHb0gME7NX1GakVvrsr+Ni/Cuh+UpVOcQQS5s7Vn3qQmOPrY12LKrc0ccXVVzEvOO
+VEq1dVZ+Na9wftqeVSXN0+uNU3wyLejmEMv6Hr06TqlsRADsfHVV3LyHJO5esI33eZD15xQhSAY
1/Fr1VZIN1NjW02/FPkl//XuVxJawr1N8GtHz9mutWqgXjkk2oIEi1HoKgB6X0877Z3JXbVNqH9a
2QOWmn6hy5mdX0Fr8x84Ocb4CQ/nojLRsSuWM0iHNEROwgTRbAXX5lYLWRtUvLXBMI5jg4l9P+GM
7wcFoJfwbzqBKNecaNARZbd5qaII2hFeGKZUl9ru2QBW0+fNS93Rp/vu9XAANqoK8bOjY6dMZwXJ
RVA/2/F4wWHYhtT2Z2gCbG/+FpwM4ywu8W8wyu4daIsngTbtX/qJ5XwUn+Y6d9PhyAbcjnsD01R7
LpvykiZQQWcS3mlzB3U39nHPXa4K/eKKVWSUJqPfWtEaGp9l08f15PSynPudEl45+BfDnEwb9c2R
WrxwKjvY5ygzHVvhYRRodS/nuFWENHJdUTuyTaV/zbmfX7Zp7shhoy+5ZvlIVSmAepuQHAz3ObbH
qQp/h6rUgPpE0dP/gNizcWELP6CUpgv/KoOjwsuQNO8H7sxN9vIYU/Di6vKcFv12dzai0Yat+JMi
Tns9rlcWdlWixgQ02floSmBgNH61Z3vIXIAsQ8OmqM1DMYgYdo7Vr/73DFRCo8fRX0EVG6foUuGP
syKcdPujeVCqmOY1HLsS2t9z54mUCXJdBg7CcHw8Y34U0Zbj+J18+YMU9F+YLsrnvXZfS+q4rI59
hMYMiEhqqofUeRYIr9N/orQ3naefoOpiX9NbGXi973PfPUZuKLa4cz5E2fANsr+1eGFKo9fie9HN
cm1mwM0REyZySzswyI7Q4OOQZzDhiEqvl0g7pmvo/m6ySXhgkD82g3/WH2IovqDqIxG4muSr9sKP
mlH1+nhpXqcssCG9Py9XQ7wDEpvXE5FETR65zulC2YtvYsCwfNh6FWoUl0ggIJJpykYW5v9KZ+Ow
bh1JYqXsu2x9fRVH0sT8Bq1TAhN4sMT2vffOopssQXmib4uQNIBKyufS79RsMST52XDrs0nPZeoi
KHkGwtxOgEfGMF9z4K8Oinw3V7pyB8oBgzT9+ZeUimpTTDhlpnXM/KshElRb+Acx1krtWHgwNB/J
LRyFTH9ilanyeMhU4eDK1TmraKn3W6d0hKGzx+iO87p9Prkbjs5bUCR5haIArTLxpXOEyBxmtp8j
RrJ8oOmQKDFdCdRq2nYQcyOta1rIsOTnIM6UUb/Bv0/4Cfo902zY2pkiVi639cnwOmLXckx0YORN
KsbS5KaTg181vEpSqnKG0ReYjVAf7ILH8gWjU/j7H3p254zoYMUAJGh6zT8X/JQq/YG8L14Ky4ro
pRTlu4cbeukFsSgWCfoxUJcW8rGdTiKDlsE82Q5ccJKz/DA4tJKEdPjfvhdZW3gJviTpKKQpG6By
l1oLnHnJKy6IXXknZebHmlWpyyX9OiZzH1Xn8Io9V5miS92ZF/9uL2pB8Y1/A4/uyxRJFxYetjuP
M9LGvzfHY5oe5j8Hf4eockY03jNIp4m0E56GE+jTfi3MZhYhgr5khPmU/Wah8K2V/f9/dRHlJ5T/
U8KaeiWijDYtyTQNI3LLIuLuZrhjmOEFKpC/C8Vrxj6D8KhUx0mz7rmX/2nVdGk2VDoy9YIGM7eh
YUQTm1DbgDtTDM/YRDdNU6BYecRzBCu7UwamAoH9IiR+vUBVDt+zsOhj77J+u9ub98rPtel9AvtH
1vCSJqY4ifrkXopZ+C2nCLD87o0vZXx2/IimBhKN2Wh0//XpbyZoIwaW9OcE1mFVr411qM0KEvC8
LFm2F80E9BlUhsvMaN6A+/q0LP+j2SAk8e7Ts92EZsGmhixH5ypMRyStjS2OzEapsnFaXnzZAlD6
JcM1RtIWfqcsdA1ywh2SZH0rovP/u80nmtyg8/XjIJkUiPUtnFppy4gri378FGRNhdVOSJSDwRh0
CLKhaGkV3diGsv5X/jpESuLOZ8sYI//GlccuBh2txlp6dDBgMDv4nQOoYtBfP0v+HdnxlZYbW4J0
niNjx5AtR3EQu/lKhUzuc+ObiaMJG/t7w5IpB+JDLq8qf7zpD6FuPDiOjfgxRuNR2DpJgLsFOCS4
Z4f/zFQXuwUi57qJqppqKheRyMSCM2AIhfF2LNfqD6X552soRxfY2a2Us/7NgX+zqBOPJtO+u7D/
ZC+TBjaDEjU+Vxi9p7tLjGOd+dwAlC81ZZ8xpBbXlBw1C0ijV55QNawUBtaWd/VrKuUnA2/uLwz9
eya6qoEaF8AS7bOJbOqKmIYIMex9brYeppLskcnoPxEP6WQLD+dMu+N6RWZueiCdqdeSYtDabWQE
2trE8N5Kq+Cr+tRNA5oSCvRtsZlJ8qpbQiKfQfBsO24vYHNKiIi5DornIpbspXH79KjwyVYCUyKR
X8quouO1StZJzt9iojZuzzgMfUPeU3Y4kPOZFUkSzUHqNPoZPniejAudWqMMhf3bEliHBYLvoXau
yYDSEAMYSffYQ7iAzxAU2nxpYyxzbsWIJ8ea8FZxTwlak0wO94QOcR8spEclm7bl8EbnqUAlyxff
tAkO8vWhrLU6q0tzcOZNV1FMULEXBW2vwWEZ8dwrpgO56BdyJLCQCvC3g8z2dqt7xoabLmhYrv6m
2vPnHlorpL2KXnPgEX/cgNN+ETGKWkTmH8597U0zfplwl+nd81bRZgN1E7b2eLHY1PHRdXa+IGEA
QgGsLM0xRhQLCb2u+eb5Xpzny5JYMd4LWrKXhmzwWiOe3N20xvxaTWVcQ4AEMTOAlfGkfWDvGv2Q
hAqnLG7rSXWa+MxHlGg6XqoTGIXvemjx//urYAcu3upndukVAiPyiJdyzEtE2doZ5tDxLaW3hM/m
PmUZXJKv2kZ2WG1FRQEQ7IsO51/Dkzvj/puY5Z5tlWFy/z94QIxh3T3DzwuKqPc7mtHUmOeM/rak
d975fXNqjNf7/Z8xws4n/iaSywY4IbU0S0v28HH7gc6XvuH1DrDYyNhMsQN2nHz2U+FUErZThRCA
7cLNWCIpXduxSMyYnwNhQ9/IqbjGU0IlAH+KcKMnaaNz21yYSHQ37MxiJEs/K4fh7FUx1QpNhftL
2fmeBiTqFTWP3vVBUCy6MZsUZsD+y4IUKJyzjz/q6+z8H1qgfWWU1Nu0rR7YZ11e0MPRyihTzOJd
77jn1rUhY+5+zAgtApjUhtbp5xHwfw9VJAkjPzJS9oeQwNesihETmJk+lC3rA3WsPNp2VBiRpfHG
Sm3Blh5e9vLz8Fm9XXAlEn6xfKbJ8YDDVr8hQjpRAeQtmANDf8FZG2uXxuRo39AaEf/w0zhqTGFx
WTbo7uENqe+m+jQiTAHE875Aj+j61Nc0tfjFoPxkHQinMnuhGSCKKoMtKsXguDdfManiOPrxvEBk
BOeVDEL1DgHotJ3vCYBDT3iwQiymhudWnG7tMOQPvTFhKeFOt1Tjn47sLXjOSMQ+jIgJTIockruN
ltpP4Uf23b2QfGfn6FWuIzso1JPixT4oZPf2AsIldGvrwnA3+Tp59jLDj54EmU54+o9WG4edmIaq
rqiIpPMwCVa8mUGXA49QTTAh+KPwP3SlZnFbfFeqxyxZp1gC7cCxANfj4otJffY+MaRaIfQWybJM
pshgymE5NQx9s7wJE/JAo8HY5ZN89pxHZ+Y4ujd0pyTbR8iRnM82pUWHhK9B14UmeLlQ57rSbTMN
YQXY+wmA2XMaGZWwx/sYeRPCZlB5Re1zTbU+x7eFYwdjvllG34lqX6Q5S+5cNOcSiXeqk01T4H0w
sN611I+qlpM4RvknmBO+4WUB0VWtlfGb/MVl7K3OP2la4K4uDLIlwk0+6vf4cDmmj3gSeDMqnNmS
3qK8vxA2cFt2OuhrDT7ARPEOkDS41yHbCoecn/5Nw1KA8rgIn4QZeFTlc4jjNl5L4Wo7AQvg2dP/
rgGZ2jq3t+Tj9XORTdJZUeTKRIPbcLajGuw5SYEtBRQpaZ3S4VKrByZDPxd3Vq7OXu7Z+rKLXAH/
rWiwF8haCLLtxXvnz9uJLqb+RPzH8gVh1FwIOXd+5Ljfr/7SEVm/vrwDatZbYtaCrrLE1CoOBdmg
XmKzexg1Vb1JkLpctYpq8pWmb/duOO3HW4oVHWc3W+FLRZit8yTj3q4CEuxXf1kaM8vEcSyRvxc1
4yhJDQzEhKFmzEODMEKswIzqWHa9kAvYi0Athesl/qxN/dTawtzQQnLTVjkRgjJRxEg8oEblXuTG
x7DOeJ4z+HHg0T9ydZctW+ZLzW7O0GCTzWSwSHfZwXDYd2Q2SBqkIzT66WFiCzO6zIXjyNzD/rPz
YSON+8VZFUW6dN2Gzvg0bbIo6XNf899E6r0gcGTltJEL2O4bVUsD2XdvM4PWh/yMZw/M9tjlhd46
3ZOn1wJ6auQQTwxWJhcQ8Hf2zn8H4Hw1xMvk2F5W8HdV3/fbuYc03v8my5UhjOEiX3Z4AjrXtSKO
18uBzOed3On4umM47q75+7vv4CXNpYD/vlrD+Yf4G38L7/ierNj0MkxbKzTNAoR3yKQKZwemd4T+
Aku5quNzq9Je0wnpZNY57Hcmj4cnpd5LOe7zG1Gi9AtdQoqmZIPtfdJGfoBxJl3Zb0cwQZSw6WdO
t4HosnkZbLcEUkv/aGO2t1Vg4BcMN/wN92MM/XJQZsnSQL8NK6WSdWKZ3T0iPXpzcq5ogWzZRCdx
IpZvYgVvy1ylS8vd5Qijyq+Nu0To4s1yUNCFkUrzoZH+3nzJuM2DjvhqHn1NXgG8XS3Z5E+51CFL
A+vf71fhkggmy3s0I9yxnB72entj3Imffs3irZUiggnW1DLDsNvOduZ5GL8d64JAMHVAFa0wRW2s
CR1hQWwE7zSrAFgKetR2Na2v4EyASnQKHevsrW53pvMDPQ6FhVYal8giqfQ+2G3OZB7QZ+lxxOf7
0NwvuWtkwbVF8iHZyJXsw8zgBqfspp+Cpl36pq+KqqvrdRDLCDaNcJHKJw7LUfOloDzZPdClzXuA
mEY2mMLqDYcFLmLJsi+5kIWBM0yRF2c8AgHNBEtwnRUVjcDcxwBO1QCkHCE/6CizuQvuGjbeYTLQ
FM9Sm0hoLdfDaUBrPG3LAZsbmYHhyz3qJgR5eAofBzQQmb6R5fvcIhykI+H8bXGzV9o6uAvDGMyj
7CxOPUxkOQGJL0VEsLW+xOi30gCa7e1mgzE0DRo6xm87udzDhtrbhrhZv5UzQiS23hLbnq2Iii5I
GY7wcjWK6CTdL+OyQigk7L8aaijtv+nF4y4j1QQTVWJhsEkfxoV8VfW/9p6naBuRjZ/fTUa/uPag
IWzDA02dLHLQ0Vs9NLD6EP2MSExIOwt+9EeByS6Hx8Ld1ggKFxCzkTXiETbwxKeQL3hasg03LJxq
Ww6TFI0rNQ4DJQxrZYq4pZdxmSSw180WDZOr7pWg5MMCfpB1UYFWCoDlAa2IzxpwCkYCZ6lmMChp
rCAkBckvQt23ZJF9nDor1IKagCJtil5vMILocIUqbSXYT0jOUX6U58/FnGo0dzwrxEZQDmMgPLqp
TP1ehSBb/+9iXMtLIVh0qDct0EflP9S/pr1QC2Q3K4c1gOzngt7+51lAkFIVGaIaFeu5vP/CzNS3
PkFzJuxQAjwYA8GB7jHPJBioBIi4Y11UAAWq5KGSjQuq/wyldhSWaaXrLVCZFbEBkqSmIeD/1nlt
iQG8VG9+VH9tdeNNWRKDhmyjxMN77AmJ4EmWr9CZYJhlhYJ7D+SZYPTIAip+NofR9mjY7rR8mrbO
emG6UYOMtegf6PQWD5obOQmCMPOxaQAJX4TNRxRzr1WTQSzchOCJOQHLEflEq3y8aRkM5+6qHZKK
4CyjxQnkZ7NOh+cHq+u89TRvbMzD7BYmTgas8VZHTXYcF9CtvDzMTnCT4AR6BMXF6SvR44yb2yT9
HPOtR6lYHOE99HTjYSPXIuv1QT43NMz3H4dq5gTnbB+chC3rx2BapNX4MptRinI0wLtHB3/7GZdd
xXupt+LOmMy8fqYUxXgdk/1FcVCcKbFBonfTyFe6FPPoud5mZBZ2GUpmW0IMvNsbNfU1TMSiWgWQ
XoEyNxKuqXCuNP2nkulEWF3GrJod8LSY0tkNXbGI/WIrLn9sDfMx0azfer3pUd1AtZXookbxyqGt
Nd01NNYVtPsoWIF81abRfwWbyJrEvQZ/z7DsKFNd5bdHkSIj8uGRdPP0J1W2nrxWq31BYD+vff34
0JKowXqwouSgx3RW+AzEiATUg3mJKUYUitcJ/C7N2VAxeYbE/PurrzjhLhocvu7RQg2vNsKX/INk
lGH1meXoH3wKUb3+4KNDGkOCrdIT/WZ8tu2ilXpG7uj9fFAhp8Ga+v5HXB+Gigap/Eg1GDnlkXJt
7AuwvSuA5lrzLWRJ1vA8qSz+OXi3kx3T9q9chScUmol1KTFJDjRr2fF85rTmuiWFezO3fMhOocNa
gT5pFSYURr/ytVVcoqdE6oZegXs85OhMveAJxAnFZm8R6H6J+v3qM2NL9OL+Am66mTE0jMjYW1Ym
+b4OfHEMUuBdOXjF7FhBVxAQwqZLJXFHiYPAoKcE0/4GBlT1D+gwM7E4xSQP8kVtVWwJg5ELqTJH
3VciINsVvaBEplV7Z4NMrmJVR0ZwtmCjRsccnx6WSu65reqhWYRgx/s05ybakix6658RjET2jPK2
52tWXEXqSv+EcPoVpQ7L+NI6MTKqtRjOsn4haJNiZaVav1mSzzibi2HU2hO2NLodXY4cCY4LG6zX
xSg34HKY4uKO2/8bdpPNl5+kL1Oyzgjdt2RDQVUfdS39hdm15aWc3ckEHAj/qv4I3FX26TgP4w2V
IFQjANHoxc7jaBJakhrSt/XXmEg0RGS7Qy+3JBrpYV1HfXOgk9ixwS67cTaFh8kAqIZAt+lIUC9u
wvDiEQ7RhvbXchZ11fo0OEwJeFrQ9Nax+QyS09tE6apnV0xFAFcN2LBiAgikfMT6ERIbiSTy4dlO
fgT+rY6gSU8OKhKgTlfceCel8UynFonjuWroSJwU1351kiFwYA3VULW76HaJg0xZT8HmpXZUaW3j
EOJJUVD1aMgnwTdneHufU5R0K8yPxWCQUZYOl/mQtZl+QV06TkFqecAkcESeVrswOqtRNagcEsRd
8BzqKwVwZoHEtGzxPcEEC9VA7jO4z0puvFks/dizDX5pLArqtF1Wzv+Cdad8bzUruIC9eKQn494t
7h1FTeKoZjbTAWE3Ma5jCqjsI4lT3G2+qCL5O9Uw1qOZxB3/qVyRx0mifQzxxT7NKcu4oq7NwNy9
9GebVBnCVj539DHYum87u4wWwwGRN+Jg2xDZROpjhEt824lxCwqtr+OBHfBf9EsPHcK5daxb4Y4M
tX9ZTEUT+ff8fbFahV+QEkI/ErYWTPJw8cTEWlrfz3heRg7pJuJjztMmgSzDT3PSaJ75DV1zfMQl
b/FBST2MurNxOMXPgGqEYYA6s/6JUOVslUMEtfG1L5EL8BsKB4bMZH6C71hSEXnZpAXccBvIWQIV
9st/DNR60M+tAQLZ9nQCRWfGOK1/1A+n83aXviiDboWEikUhk/baCt6dl7vlQrS2rz3iunaOUfnL
NiulFcPQzh9yL3by03N1Nt5SE/QIjIi4grREUD5PkRrdnlIvq2587HiJ/5MtCAaXrMENnAkG+FV2
hSKHX5ImIphJ2r7NTWCMYhb2NZ10xg03egyf8W6tdXpsT1z03PZ5ljtkqbyxBwSHzGU7YrA5umww
1CtfzT888tP85xA9CmssZbTER8+cJMFTw9KMD5iSv8vcFTbK4CfxLgVLIjOCVt/26X9cv0SEmhYN
nlfPn2cUY/6DPxZ75Li29FYJBNdpKI177xHL2hlruEfINSlLlfELUVxTGihmPeT4QGnEMKELAmCm
gVLSh1cxtZQZGHO2ULVJFMpiqDWJwuXzv6UJ90cpUybQ4kl+BSlmuB3tJgESV6/aK/jg5IfTST8n
zqRLA50XGks30IzHww60DI5Ub64qnoXs0B6Lh+LoUYQDjW9QNpVSY7DFVd53bIXNry+2829xQ/LL
ZZy2JwCKVKFlfA5AKzNKFXtaP2RMyg970DnkdoYJfEHn82JTFpqPrJrskKBI6mwJprIU4i6B4HH2
f4NOtx70zLGyRMJAUCm/BBulTJlq1wfyFOSTY/1J97pTTXIg4WBuvFHhIjGjcNwCPgHSDz++3N8I
2is9JM/VW2ASe+FzamImefud6c9yy7KrogZa3JSH2n0WuHDu+tvRRKykm4N3RKq2Jxn0BNUwpMZO
m6Vy/LcX+I0bGgbl7ewwvWI2rUZ2Mz6DMfOc1zgNVfDz7otek38Mm+Xwj1wEgjxBoyaVbS5oV69s
qBmRnEgilnpP1ckXJI13zsxC3dDrAkb12Pqy/joXHdjCj5gEVIPqbnb7XgaknB/y+Q3WzZfjZR64
gq1UumUIKh/7jvSezeAZj2hTwxEEES9RoiGa0a9Re5rc4c0C/n1c1jQ5V31szGLQVZLtrCW+rqmk
IifU7jvP63lSFYuIS9Q/MseildD9MbR5rhYYmgGx9cfdF9bjMdsX7suCXr+WM4q4j10pXT5AAscn
MW7QVFhW9acxa2Q51MMquy+DUJkchuaruaOuPxiTdrGOBIT29zRjDc3QO9fUNKkQGqmMPaUyFUT+
3w65JoHHs1BM9l8kW20UCY+e/fMNNZrsMIy9/ZExqqFPbu74nM5tsHmyPCtEx39NX8mw+hLYy4jm
NFDKgoTVlk232vgOHRsIbb6s7fmFzyXPo7VdTWGTkGNto1leN9GcJh7qBlJxZLrjoN5JaiUvtJwN
JbPLDD/E6+vcDpMBZmyerR1odNC8rEzXHJrFe0ulhuFqwUyVVPrSw9aV8OD8HCA74fZUJfT26rUB
vk5pFcoLRdaMAdadryNf2fMUatYgA6DOAW7gSNwTGeZXohOir4NQ9u6dgxcmtvFc+siTcHj/42C2
G3HYTYy6tVtrsygUATZYChMtJPrJPe5tW3HDk4utMeO3fzfMS8xwFagvBYOVMHDhfQ+RWS6wdLpx
K24durx+LfbhzickiV88bvY/JewoNmP9XOTbKFtUx0Y5xQk513exD41/LnA7cJb9NnmHOcWdYjpL
oRaK9tcQnoFcp2o/bJsY+8Iz0ry5gwbxgyb20rQYYBMTHp1XLCbgc/pfSiDz8zYPP1G1OWS30lEN
z4kHQqg7eYX8Intn0B+QwWbmi6Cy48xV/Y+jyRq0pYDndNcGYzVPCMA4UK5SrPU+kpVZHYEsU/kH
XBIuFbwQMxnK+Pfr7g4kK4BWBtSseRbvM13X6zcuZN4txmcna58XO99IpCcLV57nYS0Q8cIJjJkT
IF1s4KKVZYCR/nJnkWGLLhDRD7swPGwV+yiLRIkBO1tw0HBdTSNETcFnxZvJ3rVwhMhiTi5o1kok
egYFQSSilPZsI90V7OaBxCX9imj3HgaehNOnSodsHJP9efHSzjOwVEWu9vAsqT4rsac/yDZpY6r6
0Dtfw2NzpkFBbsV8x1lpg6mJ76k/27DKvhzGARQfck08c6gSqK7tHsdH7O563MVgczs0wPPv+y2T
LmaWjNeZsLD621KETqq+U2GMd9vBuvYCV7ym/6tlm6Jd+LgqGoj3sJCYBnVAlGSrd6GpQQU8DtTC
4IZSZqBsg8ybyjF86dQ+6IaFt/mzKoTg6Up7roBsUBrOTNRUrG8PwDLnWwQ5Zk1Es3FhvMOmNf7h
BzhyFThBfocNBwcucDsdF/D/seJeQSiDdXEho1W/7l+Q4YeMsjO8lQ2iczNxAPxkxUQwWfvys0Yu
iIudiJxFFhqBgN18si5U1hDOZfXebBfvG3gyX7Q9pfX/VaitLigWoKsRlrVvL2D3iPE46oaoN/0K
hf9xu52pu78iP0/rLwRvJFucLkOjuUTB+wBsdAs2/sb5HPtU6DnIYhhNdfxmggefBVPTNgzLW6mR
v1Y7D3apJ4BuoOE5k4RPEKKYKXkZvMig6HjRXQhQC8WPHsjCgQm1KrhKWHSwq0HSFnInTCD2uTEZ
cP3jCQ4eZkoU1AkHg9Sl8xeu50NyMt+gPXfmSgxsqKYs+Zw5Q3Q/2Y5SsOa6Y2Txecd2KXHtNHwk
5xE8QOM2pZrhH8GfbdaPDMei7x8gkKdnTXTaxh4FGy39dst/aVlEmn8lcxItrZcGJZVF5xXut0nH
P9jISubu0+2BvK9qZSG6N2WS3njUX/9Iv+u26bafuNz/jeUMO4Ryw5R0iQ+eG9hrrHZA5aYfYjsM
mxzuTmbEgOJvL0oLxbOIqYcvBci874S8YXvht7+zLtUK/YJ0g5x6S4sZKoNiCuUxJ32J3WMbLuJL
k6hEOhoN+TRuhlIPnWqN4QfkNZkYlYLSjwVDn3jxOHJ1LjJkQloo5kdWbbd+gRkFMESl4FPkz8qn
gXqBPf2VG0uDvt8ePCdemSfL5siEu53ZVcbDDwflLFrT0gNC8WInWcee8GtsyTQvdqAdxEGAh491
jUH34p4jA0oIT9hCILxLZIxkd1xBY8APpiq4lQRs88O3KXXExfjc+ePpEy+ZhS9kiZyP61isj5Kn
JlyeIzccE7qu7VCjgwdVX59aVhUS5smiBv04mqae9i04beztkcpTxUPLTeeI/2GYnsV1uno7u7Nr
uKFG4IG4z+BkKCzSqSZz1Z2I7HYauRqeoeaiKHBLspAAgcVUaQbv8KcUGvQYHpV+QDU2KKUMVJrZ
eefSdD2VnUYL+XG1s4/uKp06iZcF9fpCV5I8OrtwvjjdQMj0Kof680kbruspcQGIUp8u1JrggBKC
sL4rfJao33FMDtwwF8r3zCfJHy6/YMVJRv5k8m1Q9WvQM6UHLZnicafSxFc6MtumhSdcECEFNecv
xHEVT48npqvdauiYTSiSFy8ZoHPsJXvQJUd1bJSy5oayLSH5t6Y+9pjAICNk+Bo5ddb5nTfRrFCi
Gas7dz/s3un3f824m+6RQovQj6kns94e5K/eKLWEci8aN0yJGVy3kCfLU6/Zo359JRc8P3pSrjLb
pGO672pZclrM6KasNlBs1ie4sbCq0f8eHV4/jwzNBh9393GhyLmwhMec9yYbpD0GpR1Lyw8J51DD
sVTvh9No5w8UNutlUif5VnDZT+xhdZ/fszC73WJJz3z4MNnfj6p5XPHM//FUnt8F1mr4M4JcWdU5
MA0tXYJx2D+7LFFqBAX7Ti7MGGG6vCsSr9feCO18VCfFLnbNYDtKFLjoyGuR/qcdebiGnXWav+o2
qW76Szq0/Kt0QzBing9ryfRdgr7p4ruMx9TWvYVHsZi7Y/U0Czvs3xkCZL0dWA7XLQ9mpOUy94/o
PZWaYAAaU207VF8DjpxjyTbCISLQFJM3leu/eZvcIqVHak/sONMCRqfSucvk6uBtBbwViWiMdK/C
CTmiIpreEtZ5etTCKcWE0cptbvFnU+fh0DHWYEOumxnx96PK+id6ya7DwdcM4WfWsUl9I428UzkC
ILbEuWrEUsu6ajoexrO7UJWNo3Yc7TxW2WmcxzckRauVRq/orimjVZtyUPPXSe9T3sIQ0MGBgcYz
llePPXIkHp61TIqUrqNsVGjwVRun/ME2s7dvxohJr/WyD1k1tsrVtVG/yeXAl6zaiK+qy6QMSz4C
tDvpf3pwq2aV8WjATHJTLY8FvMWFSTwaDDwp64NMSiuGWWk1O7gbV+MHZLPCcXf51k6ng1kYi179
PzF2m14Vw+6gBUavtdnVe/l/NErKZLDH8EckcTgkiTcG1FCS+3jyTBboyW8pfJfP16iu0ws7dmUC
8396NB8bjw6dJ3qzmZW4yX7nFCX23qZCylbqKJltag1soMfeXFOQhSqtTjUfpJsI7m4o4CmHpJrh
bKxXsRBvtkfsuoLZsUTzQ9awB7bTVcU1Ztl3RZMz7ZhMJR/ZUleSShq9IR4S1a3uYnhe7TN4znik
1OvZ1Huq5TWrsKMY5uXeX5fz/X4UsC4U74uuaTD2OkDqupFYCQEOmGGaMEQ8/QnH+yM/gNC2Sukx
IXIikOdiv4TdNAiXSf47mH5+EsmVMdgxUnVPsmlhrnI6beKhxNcCVuMStvmedQ4zd4utkNRl9cj8
v49/UnpkYYftOVGVivjrutAHli4pg/SfuH7c62Jd4WXRBefBcagKBiQYwQLNSSek8jHzzdiWdXbC
JtYDpjDnaCFtZL6G3v8y8Qal1MZE4La+KElBmZ6s2PI92QP+II40vmj7HW//keDMdOCKJMR/7ebE
YKR5QdQXF9gBzRZOBB5/5nMIRKh8X2Thqxgnc9IjuNFc1Qw8umZpxUOw9JA+vLTgHwjiYTpXvl16
VDKmYseogZ9C6pC/hNahMf1nOtKP1H7pYTLyEe3RtbfAfg2KC0t2zBPblVDmyD6uLVmyZnWcfMET
JqDLV8+C5OIGWkvC91o9PlVlOJqdbEKEtr+StKgdTqbBKIZ+YSjAxzYQP85pE3JKM9sTjKUmqtCz
Gm8goObO3tIjLHl2lm1nj7EgXuIpme0AkQW+EqjAX8aqqFTZ4PRE/kht3cd8e1M382mOJYs8KTRc
TKgnoryXe+mcwzWx+aWH7Xb56+BX4tZSoq20dUykBafzup+haEnm8IYYmCFw9KkOLqufxtOoVJfF
5wWUtSURyHkHVYPH9MqeS0JTzQwb9EWBmGPDWSWNYq66MO74GeuKcGzbQp+hagsAXt1bAePQ1+hS
+jjO2PWyMN8hfx7DhkmzEdi1ifoBcgBF9gM8JPfvQIuImwozSZHsPmGy6FoUbj25lEGnQ1waVsJZ
hy4Nj6s7mPHGqHp5CIq9AZN5UgBAZb07qEzGk2KaS2XszM4zuCb+nCf0RsOn4Cl0rc0BEe3hbvWM
7S1qIjpxlDjOlLP2glyDWE27GRkIXhGByOmarXv1j+W4Cux7NRLkKPFff+W7sCWRIEflejuCnTP1
2TZIJgZFqCKPhg+rRXKW5hYH0Wd8IpPJtMzP2Z/UZ/k24AK1XzeECwN6TjwrakFYcWNZemNMIhHW
fHPCpWXE4PNpJuagnDbaqjvrCRgLGZl+wMAsom+YTXnqlBate5Z1gvkh8Tk9YOlfK34iZsnq1Njb
sD46d9dchOy2OxCGt4Gv466dTf3EEIYyVl0raRCUvM3qYHqEdj7r6v+6txbDipqSZY1srvryxLzQ
q/nd/FZ4UcKw8vQpmUGwrPk3wEB2MFCXGCGwfuOSg8RsjH0o4gPMTOckFJ1Xiwbbs0Fnw3c1zSRH
Jt06JZyN6cdodb4Lw+h87VtXD7BwHO8CP80XfEjK5QaosuYx3Sok2QOzgr/3f8cDpc9A2P1345TQ
rZpw0QGfIuUOhVvLJs0OMHu2oGcafXCfbdvK6p3pLshSnAQiF5erhkqSOVrxLyyOlx4ufw6qQYiZ
x5KGCFpwncfmUaJeOSUUce7JZtxEdeV1BY+hC/HVAPHWOH5O/6PeVSZ2bZtKwwyZ7X51dZwuRiw7
OiKZc0jEs1inE+9wLL8iDmdj0txlKhVapxCvRBoyLnoDbZ38XYyLjfkTO803eMwbAPmp/evwfKBq
P3ZaNDbxKbgACgavmZ6T+/8bFnd6nzghfstOesKD0OuZBUcFljDhLCvpiOqL83yqj9TOcshJVvR7
2tHtqonjvxy6gdDUu8fYHyGTB+xWSO6L5oAvF/NvZqcH7kMA7FS7AIhuCQow8C0AKA4hOSZQ65XF
NZSvavwDWLXVqy8xtqHqsWll08LjDZW0dzYoxVRPMbbjwycK66FPeQ2kdXptgdQVwh6f1JEEB5+C
PbUpFiI0a6BFRmcTzuH/Xu9THU9CEeGe/igonrZE94MvLYrHd1cT8gNTjTI9PEbX4RypttG7zJej
jtkTrU1RZ2JD2zhxOTJ7zbaAyf1l0plXQYYaD1M4VGt2sawLfRaq75E6iK9g8woKOcPwhw4Taek9
MgeaqvR7QRqbA4sHxXtjfdYK1Dub6ILP/mW4w6mg7b8egRgis5SWtq/i4THMnxxie6vRf71BCTuQ
JqPOgHBoqSY+eOwQNHsa4aAeVJUAqQrPHBZ5XCUboUMepMNRn8Ay6Vtd9CSob/u6UTth1Prz97ar
bX6VZsAm6Zd9tQ2YLhpLZAx+OKrhyWFwhOiueqnJsKUEmcI/mgKLcl9BrR+N4lEh0NQV1GsDkBCL
SBk8ZqDyc765EIqb1ojQc4ri7BRlAQ4QVSccNLYG8kMeqyZpec1yQzTScnVx4JsRstGvEX6Z9PFK
Mc7zfExkyczTcLY2Msr3ENmewpy7zebhfn8uy2M9g1p8+WJ2n+86gDDcBtTbuVlgaaLf8EiICknu
1Sl4drHcZSi9uHF5YuotQX5sUCS8nJOC7Z2HBUPClhc/hF9zrfMA97c3Cz7TOVbTtJDm6PmQNCr4
tt5AbVVZnwGF7zz7LI+yDdU1pK9BfLG9GXkc2VBSL4viUNxkFvM9cCyExdIBO4meu2uHdWwlQSTJ
jc5GCHc1oWgWTP2g0o5ODcMk5k77XkIZHTK0Jpk/MIursmC0vjYX7cBxQQ+BUgYm29KDiDe35Gyf
ucpNCm01Sx7ZrPC88m3EMqI1MisPD5wOrCYruSmbAyvaHlJP5UWyCCkNzFt62bB4+/4NeKuDvOLL
WX6mR3fDiaHchSV/8Xu4ZMfXaPkUmMNI3UMGi5bAZxthivAVWL3GkAotDeE/g3gocKx7CQSErKQr
oXNikPk/HRnjZV2H75yxcJNumWopRDRyEFiRQOG4kMrnJo3GcgEj/GpLw9I7+sALP+qqXgm2kRxw
YW+ohgfH/CrCOX508JNBbX0GRY/k2B9Rj3CmRBuQepmj1IygWLo56SegsaovxjT3hUNW3/oX1+V+
wo+Jf+xZZ5cVMHOE/EA8itZAIDgKg3bY6yEfRJ8BuLqkhgs2rr9mI2wBClBbr6Glbbw5k8izpZ3w
xQaZn06oCDxKftJ9Omi0mxRS7mMQgHx59ePk2GTP9GJgchApERms4C4iLpvBrKyUD/DYrpxPZSvY
hxIunNHmW6kN66y7AFOqIYUVF+NcX69ggZu0BE7fQnYaSLT1TNcVlt98H2ENMUh4R0p2CgWuqUnf
0edZm9V2+mI2OzIzvO/RCC2ED+wcEpAn+6GYXOLjatqFDTpbLozQCQNzoBoR6B58sBUi8xYAlYNq
vJ9ChhtEsQuPE5AZLVCgKRTb4y0dLW+eS2A6LhqkMqk15Sq7/OyDVmefgKOelcYI9MEKqg68Uz77
HHlUGEVvr7jv0d8U/tkVfmvggN9/8OaTaIosgxB9nW1xHUs17iclwrHaAQpJxLVD+OxbPYA5D1yH
jh/BQpkmljhq66g0SDUdkn3A97x4Ynq8rx+rxaM8/4DNP1I+AljaiWcZh9siJ+xNgkEtf4MadQh0
yO3TzEjkzfs/682EhUuA4IPZaw3k0meGAqJ3WyAl+pCUYW7m7QqgKM64ykZOBmrSK6uUgXCBkwF1
sI0IqOiPEHZMJj7IRlaK6zPLM4SkkubCLy9OzqlhvAixFJ6xvUAoFmyZVemMr7w0lYnVFES0r6tI
YymODQh1KiABYBgur3fHaQd1K5DHVcKMMWBEA3Y6TIaoEFbSnkCEy4JepyFivulVPXGBc7eXs0dE
bdj5677XvX8yWaNxaiKmTdzUEXUPiMWno4WuQWyWystfNYtepiiAmjITaUTwekDCPQQiEWaaCaIQ
xZE20UDuNCjbxeeScXUPgFNmRFPJZ/lecl7KBRTSoxjQ/qCiOCTOdIPljjPYpLyDrgHjo6rNNEN2
7gdwoJVrhMB6GOd2LKLlzVJJoIf8KxiF2qjz8WpSde/jxIdo59B1E1r3mqCnt7/JiItB8viR4WmJ
zQaB738yf05R6MrCc0BmvUttUiP02snKZdTrh4VAaX7fCwbVRJOePgbT4Mv0xj2yAvbCAbilXQi9
XNh3lJ+C4FwBcu6vTEkmXsDv7akgfSGRiBmmU4wnZuSxfWeklP9Rl6tXkqLYWd5d7IT/jBN8XJI7
dhRBbjYv+BelAZcI43ZM6eabRg+oUltkLMhyFnEbNqRJILyaxLFuj+0L/xfpQPl94Y3c2F/19BEK
W7rxHbGSTtdXl8uvh1tEN6j+c04EeXwfRKt3luwNJx1bc5/+fCQPfGAUwQKmfejFocoIOf5FNI3S
5OzVeegJtnQLgVsIKdDeTsJoEpaLEHoDCEHQaZgCv9BD73fY90HzFgbp5Lt9VWHM31xqewZ8te38
V2CcXuJGga86G/i6yvOidOVYezzU0xU5zhYvbO66D1dNkABGJcYjfvXtj4HtHb4qMMeyWIgBK6zn
pw+zC6cWBmvYqnNxuVHJra/XaWkBYeP9Hz87LrjvnIbdVptxaHqmcvkxhoMSdojBdhl76aWU0rzp
Qo77HlqxEk4HXm0kzD64dv620EydD5JH0Z34SzJRwR8Lv3MVSvUdJQCg4QEhw8rQH0Ijp0G3XjOp
fIjoV0fyE+ucGc6BGL/hfs2Ts58ZMcMon4Zg+TJvaJD3lIUZIUApOyGfzxvkFISRWBhldc74Uvnf
6Gm2eG68SWlrzo2255BWzFq8CaYUFmaeUJa1wPuICxslgDbl9xDZEJhGKXavo5OujGgP5+1kngD/
9UAEhkoDeMh+N8XoO559OKyH2fv0uVNJk9c9hy3c3hYgpXHVY+NNi9gU4BXRN+NmyQGAFaaE7zND
qiICTS10AEHl03fcx53lj6FZUsdtuNJb+XGyjcIIf3N2bTvXwPQiGAPklQ3t9LKsgqx8J/IeAyfT
3euLG/61LMLL9YHa5gw6Om11QQGyMbPfnm4NUO7SpeAqr0SwXMXDPvyN3PJoGyZDVvdP/7d/wFMv
rPJlsaCHr0ZMAWAqZ3XZWjSvtEcdJe6cU/ya7n6wHdshcyXl16H17Cp8CfYufRAoovnMdTi5+O8O
6ffcrXpuupdTG/c0IpNsaTnGl5qTuI0uJljci6ZwejJBEcLL7irPORy+fw7jEM2rUJ0UEJ3hmJlu
j5/P+C9+RJK+rtXR1UpgVBbupl1s7qBiienHh26KH+9Leg2P6c3amDKTMKS35Y8RVInYrxBt5PjZ
DVx2mNUrunGRBhBLW+WHWMlY3P7OA/ipUGb1+O2E7kcefKOjm880SgALJrjS062w27bv2hJ3Mhi2
14/fqnU7yC81ilF38o3GZqxwXz2xPizhY9WYpBrOlJHb54UEA7EMpcBlkotwz23V+9aIsxitWxmm
UWr4dK5KITIZZDd+R1qdgT/TMz1cF2sY9ArX9zD6trVjdUFqjDCPwH5qSIcW3KWqzTuoh13xcqD0
v/UaGYVkMeNYua/19A7Qamil4k0a0q0WbcLJCjX/EyNUbwR1BoZP/welebRWFitjMvcJQOYQkSXU
1EOeA0ev1xuwSofwGaHWOZo1vCbGMpKsAfNYRXsB8gpRxQUG2E+BeYTgtN6PDGgbb4M7x+xK6Am3
EK5WtWFfxbrdBdRG6Ut2kv2LirdRiGiRXVO3EeEjQgxSov3jpSctGh9vID4jKtrp+g2Mih8RC1PJ
W10F9yDCya2nHvXG8AxH41JFPFmzzQaceWxOGOEh/ewQ376gdzuaO+RnE+GYUvPI0RzMYIsK9/1R
p4mq8qmuqK2A3ZeqkQc1zgw7SLTzV98Q/V5Jm8WbZTHQouUfpwDb0Hzh8QKkYfZeJuoNY+/pLkc2
Vo6P6U0QDmqY/yLfySzN36HF0TdPY7eeJlc6QIFUwZ/95q+r244Ky0Sg34b7fhvunx+T0XMwtfjQ
RNnnJoHSvkvVuKH/ALuGk9ImRN3VC+TJHwoI83dUFPQgHG8oz6QotA4bMqbvHR5B5kLSSEiZZh+D
piVzacJZiLxXxRLvghxXvCCmXIjgJbZB+nEJ8vMac8h1nq2H/iL6zLiGw3tQl4610hpJk0qqwbF1
2KeGMOFHoiuZgYgA1luTgX6zIIHb9iW5d8j0cGvGCxsNrWApI3YV9F0e28ytXSnjS4IIqCFG86fF
n8mnfSipDUT54RUUmeoV9Yf9Eb2SfY5fhMoYiGlDof1GEGse9YVVfWdp+/DEXozWXXgwjYwun9F9
B2HJ//TpVt43OjgWmDXcxZaCZisdlbNkBsSO6AQVpdfilbyth8QjHni+4w/1f6mFgaFDRO7McjzP
3zgUOfSkX+BwBicnhxU38zeJiAfxtfToMC8gpKzGScc1MHg8gpR3kySzo6/ZdynaW9fLWXl+6DT4
6Xb36NTGg6dvLas3sI6ct1xc8rh1i8hcx8SAPLg8rZ2HeMYiI6Y5bOVus7KhUmX+zEZg9Ek/aJMw
89R1+ZkSF4DfakCXrUxZvkWfu+Pjvi+m1ttBrZwyrxmH64h73ld2GFxqEKLj7G0utsg3UfJ06/Z+
+7jydD4KaZ807iLCytKaKghmtcrKfXsFqFbK727yv/WxgJR26emSISJqWjb7XLZC68fTT5EosMjs
n+/m+dIg8r7zWSsNSxMYafTBt85dAPiNvPerAGF6P6L2c3EHMZkyyPOc9uhPV8dizfxFA/oYDqet
C5g/DNhSFHOzMmjdyMGhJpT5Gs2oNeNoigv1w3e+XX8wJhuRMOBQlcWEZRLM3ohzd1mnajFIKSKD
V2l9jDqgqKn+jhHz+brFigUjHP/voMHFZkImPFrdZQU3AgJ6xfafV8xAj/vawS+qqVaMLbBRj6u9
LgLOp/HHkURUmtLEpU9SepRy6yBoa1XfqyXPGSqfGK/0W4KNWycAxZ9MBabUAMR4xeAZZ1jGhh+k
UHOJoRoEk2v1j2bmFgMHYoqC2+mu9KE9rKTTrfKSVBAjJB1er/FbMI/Fr0QhF68jQJ+kIwwBcT34
uROTAwBjWm8KS1sPp0sPaB6dSajcJqerUmtiVCziqxdLstjRw+IBKeo2n1q08D+sTk2RqOqpUubs
9ClIH8lkajdmUaTFEniFWeIzM9r1KpQunlhnGO8I18j7llqUehQ2U5UghnRns+KOWU7VTyoi7V6W
7d9N47y/sKAHzZx3SLtdYeef3jBIUaL+d/qTNp7MNEKFVIfCk2eH6NwRmhfAm5v8lVN2Mz1YRTXi
tk9m5VHN56vKcse6fSpaIKNuMvNVYoq6APAj6RJy8jgbKKKudY6tzvM1u29QGpLW/QgM/c4CThhM
WwQR8PpQWcQuWt6kiuWOi3WQPoLNxk6r378abrT/Zl530R7a3zUPxrAdqlw9IVSLkKcZ7ggrndH+
zwq3A8rCx0OG/qHz4hMmZmya2aAtWQ458bwkqBcRutxj2zAbtYBR1w96ultFrc0P4LJpIfVDiAWs
rvudK0NQdQTFd2HTZCcjdbC9xbJ0PgaihuWJbECkfMHU/PCBD6KJ1Dle+v2f+0eaZke2qGbs8plu
PAJqUBN3t3Llt3Nasic7R4QpVW7A4MXeNw7wnIG7A3vsLExeoAgI6QEdXKIlMFZFHSAarAEr9wmh
N8slkFSoiqNpK9hIhlLsJSN/6+oKsrOkNJsPlfO+460jxDkgRIEnQGooa7CI09L2jEhgeMQn40+2
Y7Q4iQp+eFgYffuaw9gksa5ZvW1k4hfQMfJac/T4zZMBcEnkZSBOh3/EkpfkvKWaSLZMDOZSFZMV
VoHIoiG3A1btZdh44lT5C5FtYpbb0esfew0a3xg3yPrcKgsFX7AOcnYOaC3AGIZtcd5sA6ohRFCi
4RcuZrsAxSlfVNIHgIg34DVDx2ciFzF0L9y63EPqqUYF1NuZc+GQZM3bKi/XBwGP4JOV1PydyPQc
dbflWE8cXG+dUrC3YW4ZYHAIrY3tXwqUPAklY7rGy3UhPXSi9/QTI2AhcRH1rv6+52+b9hnFajZS
KWim1I/7RkwgZtY9MSSjWHCvgm8BmvGtiLOYjyJFj7F7HIuUDfWpHdUk+B2mHQwDdcaRjWtUAFf+
nqLSElia76tB0lkRSTAt6OAEbsfs+iOhRuX3OOyxUWZyHDx5CDK+7p6MrJG68/KwXimY6JkLLsR8
fu7IFf33LnMJlWAgJCQWIuX35nTTfbPNWlKeWpZU0BgMfCXsN2M21Aa0w8wnPXyE6bfoBVukvNL4
3t6zaQMAxhi7KX9IRX1KoZXqUS6X1cquu89lwa1ti8VKLK3olXgTsKBXCtr+Mzd2rkmr3WyC+Dra
lfkHfwCFjUOkNj1ZBjZRgYrA9eNT/lsf7IO9nQScBF0Kl2c6boKSiWi7XUmG78nH+woaCx4Tmw7V
A1s4a3VVmm+o73AUdKB+CrTB2mMehsfajvuPvZU5p/tuhrsk+9CbIzvCjKeVfNwRzWP8cueWQYPc
P7sNVMEpQBahlkuEhu2sO7TSFq7+yjuMBStRljQbTsT9MkzLXAOr+G8Z8B5LlyVKw4fin7SA5KxB
Enye8Rn/zJ7tcVGTxDTAfHuyfR5CsrtRpeHHG5jPa0fZ+gSZLtVV4GV2nYY9E8SlAsBZlSeYjfQi
9olf6GYvnIjmGZrqfBCuVa7X3zvavt5jx1f48SS+H0G1fPzQeESXbBysdSgoZ7b3igc/VW3q0Yk3
Uk0lbOk8qDID3plFP9QdTwrdeP7HfT0nvbr/iZO+ClQXQDEeQ5Y8jePAtHZao/HvKilY5A/qxdmV
3zm5cx7WHtOKDmN8Z6v/Y+OHN8FWfJdqg34iZv12zwEzrXzvLaxZWNrnKMAc+EJMUR4sLmSpgYmD
PBqOeP5uZoyQY+xenZ2nZgAlHCl9xq8CX2eIjRF5J0Yfr9W3LT8Lu1JmRm5+Xzth9fFCZ3pG9d2u
1Jg5Mjw5UiHbJcPX4oA+lqumigtXSf0yoHarS5Xu3sTazAtN/XdS9BCzPYK6kO6TqQFuute6jbQf
jdAUsT2hK3hLsDjT/FAVqdQrSz2GXPGoTya4fYKTpsobgluSxmJtCOyfPtz67gRQsb/DNi62+H+8
0PN93wt0e1i+uK8l12zZd7KacRMxBC5okVEtuYBXfvheIYOvuqeKEthk97Qz+F2BYMOg8Qb9CBKJ
5fV2fO0bPthfos2S0+/BLBrjIRfy8Wf3O1NDz0BM4SaULgjmbhYCmjJ8Lxhb4CgCKQjq9GSJBDVE
i1rObKewsOO4WhkK7COLZU1wdbFxyXYlAvrqfdLGI7YjvWW1yqKEZK6Rbf/anaFl06jQQNoT6wMt
lyLAdINmubyuxIHPQ2Yb+wgpDXDuEqoUhPZIVD1zZk66vP3P5yZvHZX8TL8X212cim/0skfcYiOX
EaIva66oD+tf9wrDuWcHjx1JOHb//ds0Qp9mrnr+T2ykz1EKNEe/as1aArLGthkluHVoJRKh7rMb
NLXt4lUfPdQ5nXBoY9kFUSYn83OztauPG7SNh504+idR4KPANLYiYamGu7p4ZW3v/zv6/rmMHjmh
FyypWmPddzjWnnBcUL06y6a9mmNDKRZWH80rV/Yuee6MoHf0YEsCkAVBRDl+QDES5YdU6Xzpd6yL
odML1621tSaECcL/vCvmqsLwyLAsSR/NdB0L8Tk3QBiG8Z09WzNOb0WIxRMCJx3kJPjTtjenSrzy
FVEadpyQhxl7QE+BVl3YYR7K16l/A+AJAry4wTFGWdXH46RlBc4rq53PIIQx2tAfryb//Obwn8cs
Lv2+LdsmMObAVlFdwIMR/O7dDu7L+Bf2akQAkOSdFAztMc6utfrpVcxm1pagjDbePbyU479IyQG1
BBBS+cM9nW4iDuRuyHIquW8QRNqXgA+lrJExbck0Lw4L49F60VZqDFptF/6O4i/aF+ijPs7IZzWT
zF71ucLVozuBBpc0bFqevL0I3+NGad7kn9XZaZ+/A2pv4QVjOF4j4XY+TLtb1n22MsNbHxyyN/KZ
4JvuSeXo7mrlu0/P1cVX6KskjnGpZevuK2MVx23tlkUYJNivWe+BZ42eVBiOUxeF5rFRtMenIm8y
1hP+R/qAxFs4k/SgvE7UqcC6w6FX9PjHxwBsGkawpxPNxKFeYPGSsUPgPUnVFdjiGKQgTicaDhSR
xiGkjdJbQfHb9xf1QvgOR1SdtbIt9rSboHsRF0f5KQbS/r0QPslTMUXepbfDI1AnZrzzTIPOkbFF
V01tUUr1/Qgn9Qsh2LHVQo2Jgf/JGmTAI6P1Z7UZ3c2Uiva25pg1dYxEtDkvGE3IV0SrRDoWXPRa
uhfcIutHBrFNBj/kMLedaIxys9xg5ikzee9vi4sBsrkyW8fIn3AkDD6vAcB+VYUWTMUbDA7mljpo
1YYb7wUrPS8AWaW9Hj1mn87ie+UwJOcU3d72Zx+QuDOKZFdIlzdPVhtF3RWfft+pjFAf2Tt9DvU4
npRb0sdqCJwmE9CibcxdhVyHVc95ILcmh1slpNndpP0CQKXcqrKbHUARr9JVOM+V2lBUylhbYY2c
jUeV9Q250gWGD9sbkp6FP2tUbG9NIlC7FE12+umQoUSS3v8P7qNKTKtVz88QpzBl76A+sH5T4yso
hQiWe/ojdSwKGYgNF14YeM1wzWU+Kvskg6Rs47Z5NQEAiWg/uNwk7O67Myl2nIc7rSmQISitNEhA
JvQgaca1r2n0P3MbAc7S66x6lsfx/UGIXaaZoHSIDjiIfmV7/2XvaK+0SWggsRKiADIWwI3qLbD/
oiRQjXKnUFUC+KhmroK2rnkEvS/HQVercxIswdgefD60tvFUiCLToaoqVjF6WoCRm0QkyBu1Iz1T
70ZVrVUbAJUCsFuFeD8lhHnF+lanA85BCIC+6LyxV7TQeLPtAHQ1jq5uaZlvV/oP27iRC7va1htQ
/e0OMU+kR7H/s7emJYP598dxjMcV4TEP7dxLa6LAVTr0l/m4UE4AKlE0rNVYzNambATfrLKn7a2k
8Foj87aBfEBkBbMjFgPPQobrpCYnEw0xXfXQXz7sxbY8MCBb2DG6GjEGy1tjNSqzNKS/4FIYzaeI
iLIYSwhbOiKXRrq9lSDk5DieNAaMBGQ/Y2zwxaichs1zuWUSUxvQVcP9hif1Xlq/h2D5jZhnrqzj
BbWSMd8rxTAXrBhsaoVIbjTcdiW3wtEBUEhAnjFIcNobT7S3hSpGsX9b4ko6+RL+HZSsDAXQ4fT9
IjQC1v6xI9y0qoxAauZfEFnzJr+jxwwa0STxXAej6KRGjBkQSlhoVCOw1FbfQx4zAqqzUGxnmdSf
rW0vNLmSPCB6eolX/zfI6WSswMIg5oexDj7se38Yegho5jIOLqc5cdEbUXbn56NYWYM+qoGG5NLC
gTAtvACq/8TGni3QjIBgudMMbWWxFIOUrrOVqFntj7rBzpWI/v+zxtuTTkO3dhgNf0YLQfdG6Tgz
nByF/Gp9a7nj4UilXin0pv6WY+hZ+N+8Eisf8YGo+QyE7+rbicKySJG0WjX0pV/ctUwpjhq3vT3q
AozP/xt5F+vCyjAClOAsAXPakiGe1aNqkkTvGGNH+70B6Ol3Xpn1u4xHeEoRCI0Xx/g/GjppDdRn
1C2Ic6hDSmhNa5IFW9xty4p3+6VpLuwlfjnyn98LSeMtOvsFyJdsN6ddRkX/kLEkVZZGJfHZafAJ
+WzTs22h7OjSRxHtWRLnI0chw6yWt+shDipq6YrVd11Wl//QRW2xNMDjAs1KYNKVvsN8U9IhpoQ6
EALfBU5FLaRoery0KWyFYgIGYCotfBspTrh4qET5IVLT1rRsTdTIfMC5DKPIo0+iOoyhfvuZRLqJ
Z7ro11r4oQZqS1VM1vOm40jtEGszWuFIopOzsNhH4p1hUmeySYWlNXPSTF9WhkRQ/Y2lR0AJLWWW
dSAEVUh/yLjAtrhCIQcWxMXJgm7/5y9nmaDgkI3FqmC96r42GjEvff+RSkc8ulsSVqdabqIviVCS
OQH7kNrTPPGCnb06wBInligux0q2Nv4CnbEXJzxWWNMhohlqTKWcm4zMIIoZGPpwQ5AiVY9IxaaL
azYOdjOCtv0ynIFilghi/8U6RGatTaBMZe/mKKSma6oGNNHbooCFdRH7/9YZhdyx227j4uxktcW1
sIimXUQo26IcBd2BDY9VY2yakS5xkvKuZH0jIZrfJf2D2stX4AMUjEDc4ps/FSYmozbFhaCZSWUS
uTHaqx+lB6Fak/ehSEdMaXQ2pVIFXzmV+vJvdhJZ1p45eYJ+9CkUx7owrd5KGRIAs65ihdc57BVv
ePfavN9o1zWECT1TMDzGFOSWDyMav5FTCvB10k2XdElBhlbJaY+yqm33oWe+Brm8Tbyf5Zto0KGt
Mx8CTIob+ICrqkW7yzQIlpjllrJvWQ5u8WHpMzHAKy6d/sRHNgAv7iNJNmDcEL9XZi3wBkd4Uxli
WrMYUURxYi5wYb0ua8rN8W3Y8gVrk3N7eoXXhrzfEPFV7EpYbJWH9ryDsE7e1PP2c0gS65FzdCMM
O8TLoFw1grozSwh1NDvdLVxb/ZibTdENU1Z47vUMqJq1U51yam9RG+UU+BdaR96PulkZwydTP7mQ
5UKk4mN3jDTRXvDrqf/TQe8GHCfN6jiBFpUhl+ouGE0H30GdJMiqphyY7fcYbMnKC4mWddOfQljW
0xIjtvRucOUtyTrV9xM3wMhkl/mZHszR31aYXwJyZGE1pFNeeJCMw365+J9ifxKOmxop5TJENlcB
IFDHqkJyhyzO6JoA7hcEUlk+HkYsE+Q5A8pBc/0XvVUopxdcVQIv1X1EXF/IaoHmaUgjyoNRzA91
tfAJOqHKvj6Gm9rqjwUPvbQ3hKvhW58TQ6UBxN9/p1nXYlSEj6COJ375TA/nW8C0hq8+Ldr283t0
IbLFBLz+wD8xbOx+0dRmjLb12mB3h5eGbYWrzzzLopd8n1ROX7RFE4WrVZNJ0aFhAIgeewagAyGc
g0pd67E53iY797g+3VTNX0TyQk+X5f0GCSd4RFg0WJF66D8VWPQ2pkWjC0/Ue1IvylMBvI4m/frw
209lAOT7VLZx2sGwic7RLdkzVj2xyxlyPeVt6eULR5XXPdfzoJas6Utbzevfew/5VavUe/3lR0fY
xy2wnxxMkVCmzJOaXOXl7tJgXdnte9Jc4L05qDmJCwqJUNPkr3Obqq/lWI8fD8q6Tq0TY9O5J/p8
qoT9glgRhIFsftX44gZ/Dg3cuLNuGTkKFQXvgDLzJwd+jCnlVHLhw4XQjbYB11ZGUjOJ9bPQxVxQ
dKAdtx/cdAylKlpVHzcvKkq7Q0OB48LveEM8sESLrGUlPLl2iXt4ibLrgXiv47BD2INCX97CaQV2
iAzfLaqtj7z9Mn+jAtRcLkCce8X6em3AZXyMysijleyBiWPzQp5Vk4LVD12KU6RZK3g/0aV0AjAi
cKBpNg6Xty/2+UVhQS/lbxubGsISFhmgaYxYhamQGILKa3Cn/c9vHVD8chgngirEYlw6tB8xeDfQ
WcMzKJHtUAv6KU7omQuBrT+kuwO39MY152SL4zBY+hgi/524GAmK/lNhdMqkyzTypIEP73HFMVTa
81jO7Y8j6WOg1+YVcgtjUwcAXDxanllOheZclQ9TQ7WdIbqNcbAYtgT/nkNA9hAJaT54e38KYj87
yaK0JUfUa4HqcE1oCjFob8jg9meVdooY5vBrR7W1hOFOWc+GPeyO0K4T7JRZThrO1+cx1cqDSI9C
h/dyJCCBqPi5cuTF7BnrTcFbwXZSaJNG5lSH47EAm7OfX+TOEsJ97rnKiHhWffkcerjoYtnVuFks
1Y0zc0cFTB3N1uqlIyEPByhK2RXDjcSuuwjSF22wBxKEFRjEtCqxXFFAWqt2vz7/15uhkvVa8HYu
c7KA1zvhAHBdZevyeB6iFnOAooQT5ShmAcP487PcKbnwTRBi1pamBmx5/Hr8HEcN/KbWt3kC6n9S
g1kwr3DbSCAEPCDCaGwj4br33y67bz76jHMeoIuco6jKbWfRqn2R6OsEnaEH8qdE20vcNwXRfp+G
rvWghMRIUJ4APHul6A9+LYyRVSMwcHHncuq030sgSrbwOUHj4PZrYT8OAYNRvQI84jW6ZJ3dea/A
ys8XVzUUvGmN/wpme3rICRz742rBZkjNHOENfMQ+7ymFjGy80pI7OXC1txCYNHWHrmYqEF0lK+oF
94VMlIgqfgpKlG6GRf8ZX7+XQdhNKeeTzge3pn9XnJcKr0f7xmlToFCTpEZMVNnDygstFfEoOLXW
AZ+NwF03MQY3/LZ8elHRzyMvuqFy4zrHHM+Bo6IwzOv9XXY2DzBJrYOVJDthhileZZmaNRcl2jAr
SHmo1MJchVT8iWqNgmzewCn+8vURpO/pEPPPuoev730bM12ky3WtaclUuD0Hbw5U7euL40QEfu5T
o5+P+iZTi7wR0DWQfL4SbNF4UtsMwZqqTE0jRZGjLVCSu0/cAb5912TFNhwtthcUnixVUb+hgcvl
bsW+Fqv1FRPyQ7FaPthiR2QZgyODC2bk3ukSbp2O7Ot2C05FpwcQWZfJVunBgDyVQLNbli2Tlxs3
ne0O+cj4KFaQ0ZvJvfnuhmi8yknJKyU3Z9mZR6IF1TCMO0zi8mUGaPmqoAb0BnbSKFHf0Fjbkh8S
UWSRIgsLcOcl3bhAqG43nvVxaeDfInhAEa7LhLAgcOW+U6ERWT80rvFn72iZinCzFW/t12+nEhhF
+0zC3WFQbNUduevBhJ/lq6xEqTvFDYZ1SO7iUvYQ9ukeyanA3M5wfyhQZhUw3unzTWFFeSfQ5h5y
afTQwVt9IiIYOzw58PVuzDZmQ9hB+DjcyLk3o5ViAix1LqvZpUXAvk6FtZ/BP1JFrtWCq0LgenQj
9xo/B85i2rppkfpGrN8hY4ppwmMR8fse7aOIBQVwNp6X5iZ22s5acWgeGU1PoqJtiJaHgHGFYSgf
LBnGz6O+Zm99pOuzy0iHRUuqB+3Y8GahsHwZawI9ezXnrxJ24B+3sZqkuK/cMcddyMYF30tDkqkR
sRrBRzXmHAEri1SvKhrE0f5/6AE6HK/k9OVOo7+LwcayxvBOKlNzZvCtzyIzBrLaClpRnVTPyjh2
My+KEiP50B3yV9I+ciW//MaBYnydeXSR9h03koKqJSDDkZnlE3Ew4VyfI+oYqbLGDgoxJunC4PVW
4xQANoniKtzxYXwg3BsmZa+St4Tgmvy2PQosUI6ax384iGvNRLUVrXpMbadRg32gXXGCN+L5JypI
W4SOhBoiNCChhL7tmaQkQZnJ5JXEYlysAk44rx6wki+o5M8J25IfmZ6SgFnSkxuS63JXAWn/wDYe
EJFPlCH8V2CtIa8Vq7zuOvSDu262txm72btOfgU0RTNeYHh/0Jgfio2wwuPxGFNc4WfCcS1Q3Yyl
MyK2nTzKpjmF/wsD8W0Xe/LdO+m28DRSf1+RSAkBiVXh8glmzIrXj+ORJE54Vq4x6O5SBf4zVRWI
XKhBiADd1ijkyl9j2v/BWwfyxu2qVGPY0pV9ngnZFlHLspHlWx+y3vCsdMaKwsWkS0hfHG07058q
hGDFXC8n9I+Ibr6QdPyqgtQ6SxvMlsnt5H/dgAr4XDCVv1ddq95bpmjrwz680The2R4/JpQWRPJs
2FLRasdOQJ8LR14kiFg8VR9ClwiMeS69Fw+vA9Z8oHm9Mkw6SRXVdJEgw1VyGHuUwS9Sa0e324zV
kuM2Bm2GrcJgYk0gwxujTsf2lf+rGJvqYXq/bU5Uak3xLack3Ylmq+Uc/GBphe8vRiCcyiuWaH6W
C8VlmEQy9Q3w6Kn/JfsPCsBHhsDRrJowCMWvTBgFaIOezvW0ecc6N4RhR2viXG+mR5pkBsBJULM7
aqYLXhCmKgO3Mw7+K8cokU1Mg1DymeTN6rU2jBuw8txEDKpkcwml1PHkJiwOr53cPE31WkCwmdnG
ZLg/8oFa+NaWf4jpNVE/6dOILyVN5ITDK3tAj4pXBb1oMurcGAhbKG199sxhOr8WV4lvAFVwzZja
iV0iwPLXA0KiU9c5MBScvrmUiC8venpRRtEmmNoW5U+SlorSSSkopua5MfBvJ1pQxJQxu4BD4sFc
EIWYLH3/G5E38ryqS0l7Yy8wIiWnV+ndAEgVip2GKKDaYp6zWmbKpskBkbse3u25IHA/K4RfISDh
kVhiYsiPgR6AkPOkTRVRdxXLV2Rr3O2icCe1Ktj3l0P1q649/8rgwlWLVH/SmV1lBR0vq2CE7fpv
0OCKZO/ELd+LtjYgkUt8XAzSB5UkOpgpj4VH46BJTdps41iu+nP+jwOCMM+/dbaDh4mxIDn+gs31
tszzUQTeYiDpgQtBKsoXH/N46c0Q0MYDExd5A1szo1oSkBG1VoAJlF27cP6C6VgVd4gMtVNSl5vB
3J2gNkQN1lSX/NGzSnCgEQ0FZusH9JrK/kym0tXPSOwF2MNilFr0ykcHhvtEZ1zeisg5Ew69VU/R
hfJJ3Up+q2uibRM1g7euGQcPUdOxAJo9J6u/SDeqzH0nGBgsZCbxjGZwzMbHhD+GpC91kSWouEXJ
/g0+MtnTKUsvMvrcwGulA+uEL87ySZBdalTEJCa2pTHTZjRmyJkgKu3sbcI9xnquyq7cw+eXTGYf
saL0617HKWdnerVywCpsm90PKC8ixP9/zwtJhQp8IbaSFfq7zmGlGIdTfQnqFCpinv/5wmtJZ3pP
bHAlX6d9xZPNDuafoNX7AvDMGbMBYjy94vWAJZY0yj94ol6ohFEn6Ho+qYwRIgj9WlsjfPwbTiI1
clwKimxFoOk9FOHTO1Kz7i74YX6GlM6L3QxpGf9aooH6R/tZTCbQE2eGWTc2njgsoL40TYCL12BR
To8Z9YKdAVFRCYmapRaxrv19zpDVbZW9wyFYma5iY0X3g154a+LMJLvNCvcNt2FLTq1iuZNrp7QL
QutL7PZeCFX/uwKjJQZ+S6dEtz+x88FkzGtIFeY2MLNm+WVWa43qD6fPi0txYG/CaVoM81CYC3Qg
FtuuSNsVBQIGkNsOsVgNrejUOaAxtAdpuuV6wzI2vfoRztDb3jnMFUi7V3ECwzgHPY8JwG7y16Zp
dhCFhJ7/Wol4U3GcpCgysszqD6J9ZDWoZXs8Ya1v4TVj3UH33vvSkrKCRLlH8n+DbUEdKemQlLkE
Lqw1C7STcZ3HFJZrr3oe8tDcDENP4Bn+UOb2d+dollx9XwMrmBR2/5bThaNskj/eLH7a7tTDFFL1
DUv4VB/129ivNOj8k1RwIv09XVLbCUKeyA3IkdtOs/vj7KQj8K8kRNtBmjwbvp+gZ8BWgGf4+iBG
BQjxOlbUclLONPnINOP6qS+3RzJo1bzeSNY1dN0gZd45n07jc+73mlIC6p/SLyq5nyIMFnkkX+WQ
INx3VWezNfy6VUUvQZPHnS56h/rGNLA9hazA455Go9kjlYihXS57z4xqngEikxzVdfFjHo7kUuVG
bUTBD5EGY+e8WaX04udhcm0sl8iT/iXS9F/6Mvclzbq0fx/9//ndTWFzUpPWChnKODWp+kYq40xX
RPW4Ey6nNjnxisSafQpoKst0Q5IVXFMXxLROMl6/8bT6Hul3625tIg25Sjy0nhCVAogiRLE/Ohvs
BZqxLzVefAh8pb7Lqol8qehPDcm+7OgZDJCvqkYMLG3QyYMcxSfHC4hRDmmRmYIyl6Ua1fPt7O6S
p5ZH+zn94cVfD4fgh1U++TTSKi2Ov4N4mpVGVoOZg9lVJ0u7IWPFrRl8RihTKxu77ZhyvYLn4YbK
Zcx7UdIuhOYUCvlHpsOgJhPNTLULxBIU/XheNrVGxxGxp5hlTqHWoyWZpj+XwNNZJp5XCb+u3R5w
KfAMif7OICsGGvBV4GIlbZe2lukfpBge1dM0+fwDeNIzwc27/FtxxvmVfStD0miiPqU25qCCvLVp
xwGgHSb13Q6ro46lzR6zmQr6itGLyt4WS/t2RM+au+9pn7SimMUZyxynkcJSMeolybRR8hYxRklU
ALOrW2YdxsXOSP6Hfu759h+oEZ41KemAQej0mKt6Eq7gUhwDSQ5CHdjfQ4RD6tQns5x5+fLIEhUR
8GgMSVUmx6LmJm8WB57cRDxWuitF9C1wn8JgQ8FFjWZvcpOKXtHBPnJarSzqVl23V7fRZDOaKw40
D7Jr6pa+j+Mk0InPpZW3QuzIfq0YPJM0bcfemE4m9Gre1UftHpunjNC8xS56H68VZoxkOV3uZDkP
lfU6JrOQjgnlOXGjEV759BaaooxUDJmLkIPOQ9MiZCLyL6vclwcux0OPDQRreaKHNZzGpAPmU+cD
Csdc7om65CMjRxtobMx7YBU0ub8S+re1KPwMQSwnUec7HPTL5VyCzJHFhn29BdKFdhJd1k9kLgWu
vbrBhaE+hjAwbpMfzwtDpKjBh23YQil4rMpweeWY/C5+mTmBBKTlrjiHF7M8SbDZjt8JpMZZIGZz
TT6TPGryfr1Dz2NQqoMwpTNbmJ/ZhWAjrrcWb1Pr8OR1stYPAfGhXoeccqB0oZZHC2dfH1Z58fl8
XlKh2b3qN0UUo1C0X4HL/pZqAcSAA9m4BeFDcqdQ0UmaSMJ02GzbxjemM4Kiyyuj3UM4PdncIh+x
8+eBxrnTWDndknTulNM1FC1B82tBDs+XgHVHoZR4PflC0Tg97lNKmmiD2zOHczODzeNu0Y5CEO1e
HTBsQ1Fo/O6qWRzG9kfAhbHtHMuV6Wzw9rMXn907G5msK+mllBG1c0GCTgUB5mzY9dZQZJy0+uI2
8NGO69noHIL6HGpc9XgEiEDNxzKp03bsJ1SRRZjkMegWb50RzutZtZ+kVirD6rWj84CwXxUVlGnp
tTPFqNPOkqR4NvZZr9B72kqhrdCd/BO/CW9ie1/3HTy0gGJz8Odo+6PSpWiIyor9X3aV4EpPvrJD
EjX/AD6jWo3SJkqxPF9v5iFSXK9uZTsLTfzx39fwwDatGcfyomQasdSvCamZm+oLqAZubwJK9uGf
ryfjcIHPrTAbf48Sx7YQ3OBrqYrCmId8LhmieA7l7i4rUh9i96IEcShdSAu9ncqJ40HjAMIbSGu/
xIRFVu3+7nK0pjvlTyuTAULeS4H7+D1jUgU8QGBJpGcaJn50oUtdaa59Vz5bT1cA1CwaYJ24weov
ZGt3Gq8cpsREbfQYFIwBTfZzOhtd+3wXfQmC+QSHASdQXRWmJOHvs0WhH/bDrMJ2H93J8pFdBScl
HDTLPC+ljeMjrWtRgmZTbLw0jGGWxdM9GocHOuvkD8T4fk5OrBo2KbBeRwLVXCIhd6zg3pl3HPac
c0q0w98mkWLL+Lu6JbszRQdQoK/GjiaAkkAYfTejBRBjBEWdl0t7DAjU1gKFSANuaZqUVzXdcD5N
B1wHrnPN8XkB8uXsOnvRS/SA/VBwt0cVgzb/L+2qswRwJZJaB1EwUoVxUXgdHLvKV0QlzlOi13hy
AdaUx7BquaGc+DNATAbu6CDdlorpb03EgAygui9ifKaSfMHh19742l5tDMzDAJjJPANctYWCckVl
ubusJ68pwqZNIkjucFOJL51SjpCN7wPcO4S9yT5bPKg84ObnwQ6757/b9rZxhTmDZByX6tnDytI+
sgUwTVfx9MJ+fDd3RJLFURHC9zHTyBZDrj4MFfeOfR0wc/KQoibImlRgakz233UQy9USmPOuXgUY
H47hB7DxqZSBuKlJuJpSvBaMeIUCpLjmxROFdJO1PvYkiADlAQ+u6dUZARrzhGqY/0NJTcJvaQ0m
RAx9S2Z9TnUptCab8xgs0J07zXxmzd8oXcvJWJkS+E6M1vWsHpMflqCnXrraHxVphczRbaJjKmXi
BKzlGxrTaZd93JMJWUGRqY36mx2wU1aGvoHTY+k5MhRcGrTRpk0oaiaTfTYFBnbZ/1k+xlJeT4TL
fxermw3Jum2AZS6PBny/berC3RJtHSqZfq7PxULm8g0wtdhldlkuerG54L/fpJ8Mc8E07EEUt88o
4qQLafQUx7d8xzJ5Ogtw7bY5jTHkf1C736rQ6oliKEj2YXS52TTfd7LdD0T6iZsYLCXF4hui0b7G
IUAubvwONFwughBUKBRCmI61jijryyWTsXJMI2ziHWhTjIQFColDlEIISE7fU70N2gE+eD9qqgp0
kLYCjh2fQaJFB29uL65ejADjDKBs1gCKPX25iFw2HKgUCRxzk/yAdkdXeb2mKnwEWKCcCzfSOA6E
pPpvGQPAwKfkx+fg3yPXLtZPzIe02pgULsOE9UoOWJL3X9M0Oajq4VwSQRVdDbdtvQBZhvTxKoO+
+IYvQ2jtOytBDieWohJhmZChCcT75xqsYgQDFCUOwK/wy8fALRXeZD8aAQZQYX4Tgc9svlc3BnjD
7ad630EDrI15NSeJvnGefrGz7NeO1FmTt+nr2cA2dyGsACiSLBZhfPIdxCj5mtmzFcMkzcBjwh93
YBclZnvorKZHkwHNpxJmjUkUrxBC9dwU8D4PvMCGGNpEnuBw7Z7U5GC9nQrzNAE1gTSVB+uQcyhX
3zs1/yl4X88i19lw4TeIhG99+Fvv8KpMbZF9RQOBNp5L8rkMkEY9nLZSl59BD38Kk+si4O/P33x9
d05HSTsP1gbBJ8/x45rD2wB3L0fMoxsNvbInvCgISYYmUD+0UPyKPeeGdMO28eBy5fTf4pPTGubf
1omgjnXDHWx/5bxT/DJ4g1bXSIWcu5pnALXY4hYvNbT4zIkpkm0pLvVOkxrZBj+WQbZxFA8edT1g
cA9v5gmGegDD1aplCOp6SfCt1W9bAqmmInorXgqhUv6Hc5B914onYRkUPzPXhw30cNlUUCLC2kGx
dDWmRxHyQZ5TqsbLYtcVaegK7y1PtF75cSDLNNGk6fBhdpYBjcOw4xdp7eSoQQ+o+cQWd9MzQCRN
v0NWvbsw/HgEl5Qj/VhyPwylxAGTm0Y+LXvo9w9HBx4H+zs0EuSLEtoUgLDweu14NISKeAZUCA9b
Rkty8A8hNdW7KCbm7utPQRFZHpy/P7nAGVJyhXB8fJI9Vfrv3Nq6r/k1vEakfFCHJiIJOPlvfgd7
q9lf1zhKF5UWR5eIFH9MJn1wV7ZbUJ7ye9euoh2MaLkOMzc5CmfSDH05+sbfIS49gMupmbNaEEgN
U9TSLiGxikjv8zZt5kmq3ofFg+ZNzE9rs/tx0yfOrpyK6v4PwuUcIALT7v9ihl9lGBfxoYM/pU15
lfxaxUVTQfV+cLEf9jSW0eAz+o0nDHjjNxLdVb1MrnltG6jurkt2MUxhAiajzVmF+bmadH6M6AsE
GsYAJoqpognFdXMgR9iFJpRex2Wnw9Y21P/MhQNnsSkx6hgZp3pXFAqIIf6zOOmIlPTGtDVMScYe
0uS4ctyvHTsC3CAzt67sALHtHYWa55ABoZU/GXVnHNjD2Uau3Ldc05sZv0Jwoo4mjRCwf+Ozbrhz
k2BtideXfQaVfQsHJ4UaUE97Zhbfkc7dK92hZNVgls9yx+rjKfepp8X8aFAwpHFk8keJnw9URT4l
l9dbH0dBfU+FsRpGb4+fqPWUwislC2K11RiaH7oo35Zkuy0t1cbGwlYl0nOYVxbwvtDDRQWmLgF5
3rP+Lcrj2JDcr6BjCmpIIhbch70cCGsdbFTJFZtumL2xYDdye478Ez5QxhJ2dckkxdFRjwoGlBKz
ztwJ3F1mpvja6qFHqBYiNlVOoWm//BQDMD26xQK1tHahNnKKMaA/dI7h+ivg4zZkek6TG/uYDs6/
dCl4VMcIumZ5EzZ0LujTBKITXaEaxE78WST+8tLIWbTlRvz9D33PgsHP2lLOz7sihg3cAVtpyPMb
Y0db0Cl+xNs02MhLcyHxgTdzlRia4Vy1IAsNV4lNrarrWUln0MgTnHNL6/96abQgKrcYipKjfx39
2fi8nKY6OmzseGc1ijl4Kd6AgpZcLLBZI4ks+NLDebE6xFhDVwMfb5IwJJmRRePMq4O4PjVi4SVq
M1cFcy9v1G2llgyn3e5fw7kfL9VJp/MZB7tbyXKKzHF0Pk8bo3v48EA27agWLHiW0Bwm2I07IGLC
8qYNXcqHdP/dSay/hM/osUAiDAazj/BALtIsVDow+ZLOi5S1SPAovZZa0xsD8inMzk/IfF3hRx5K
PYGqFRA9BvhGfFebp4uBSDDYxHa3UlGqOpQrwn53LgkTtKg4POiSmrXmxrdQ2cych8fCxsMQx5r9
g+tG8Of1iuNeNxvzJGxW37jk3N/gJY2P7N0xqR4DmX+WjflVP5Y6LXfM1A7ljyhzYxJy565SZoBT
HKCJbYRmoIi4f7/WX4W3aDiFKzzNnXHCLX7iNAUb818rl3LzQjz8dEApGpfzLat/dx2kqFwA96Xg
4oXYhRcyWgEx5RuXTVzyc68tWntVLrF3Bl93/NcZNl5vxq43pc4zDHE2CtDSyJ/2jHUvFPo6e6wM
OgSJ5TsOn0FN7H4qLtBuw3MuCQ2zJ1HcMyQSnDaas7Pbc/y1OP58scUnguj/rWk7I3Kb5Bu/fa5w
njpY2iXI5TnR2EIWonv7LnZeaQkjeoXyCsN6y113VGffaj0dJb4jy/VUhJ2wI3MHeU2jEQTezx5U
X76As3iwyCr8kc018KvehjyAFQBohTBddxOkhGnBlvXHOBEl1zjbxWNdzykg2I1vavn9DX7Tajl8
hny3crSq570xCNoU5XtVYwZJh2lRvcdYg3OO51++E4AGVfPCZIwefu8A09natgG9w8DUW3y7o4qn
L9DlrpvMOr/cAZavaj9Getx14ZX53NupsnxNrQ4BK29mJJYCrDVd6ZyWlH30XB8xR5Tx8m7NM8pQ
fMKbD4OKDJVO48kOzfmlW3jVOFL5DSzrihQAyt8QIGMKQ0WHuoklk4ox+/tWyKeC+Sz20MCsEQ+Z
1cOIQWxJdhqm5zzt4LZyU++cXXyT6sJLDW4EmNy2hqkdMps8Z2fuc3jriNqzvN8y2fgbDVJb4p5F
yPG8vRVE2cCx47W5SDQPQRlnUYR/iVwGj+fD6WECHkr+lZlECUEKEEnteQ1qp4CX3LEmhuSf+9ja
jk2nFg0DFez/xMiImehvsH8CXjiByQpAfzUtYn1HelyCF0r5ovJSFsusn6iI3YIh5UGCefiPTj+1
M4G6tDr3y+ZGuJoTwPmoGT0M4chQv56M8R+FiZydtxtBkiOWHNuKx6HOT+O0sTI6I7iZBc8/3iZ5
qJHSTHsGPgAgZAP5KVXfqxHVHZz5oa6JtfZTty++gBInogWPljBZB4kb48a0Onoa6Tpt15vpggZn
ohnt/1SlH4fUHxga2cj3/1ReuRRs5DP2J53U72dePQbNBA1hiTPO1AokA0Pt7LcRSmfo+KbOB9Ro
QPVsrY9AqBbLU7C9TRnZOO6K2BOQMoo3pXIuPPG/xdGV5HYQsjSW/D6lb5WAmwwYyiFAtYEMFXpk
QrFZgvel9dGhi/thPV20nWNStK4wZ1Mw797PTzcK52izpv3N13X2pnPxUygwujt9Xpd1epOTSimi
c3tUFKDcbTT9qP9ZinyrW41f4r+rmhSa54m7xOmnnOzjvujgmMGDLX8l9Zo5/CysXuGkdtdmd+Ut
L8UUXid8lPhU/I1JHDBm73cDWYt8tb15LPSjxWKDRfZp6U14RPYp9MnJUoqSjS0zq69ybvVaYSmR
lsPL+uBG9nLv4oZWQZvzRK0CHWro6FCMu2yJj/HiFtF1XxF2Iucgo9DhLd1fZaDbZg/n72Y9C48+
1prog9XveRC8I2N7ml1CDF6iUyufjNbfretdA5IFJz5GmF8nP4l+vzLfuhl+XGc8CWAOYhaq/m4D
q3b1fHoEhoj6bldL36vJiY/YN+KoWO078mE9C7Vk9zTtpYwlZy+wYYF1ZW/f/j72nx7dmYfHB4km
THyjFfC3OBCyYZU8Z9zoOXoF6MOTScpONHSBOmZQOEziUPsZpLW4yD28B8Udk2EpKeFm+8bBiniw
B7/B1fZB+bPiSKpbjhXXpiBFVguX6jNrm5FMNSJRHdyj+P9Z+zEitZcyPYIOFymFaGz/SExdMNkK
NVYG67c+D65hh45r6rdXN09gNX9sepf0AxEfPmiNmkDqRMGk2Ai1fcMTKFt4hB4EHa1+Jx6PfR6D
iEcIP3tYm9iIs6/sao6c7wbABautj/vD7LHAnM/ms8KZ2tIJG/VVKjJsWzF3NQctgxlFHAh+n9eb
zVKQtziDoeSx/N0F5TC1n2Igo8js+z6I5uSQf9kpgZ0ie9BRZXin8YeRK0mYTkmb7TRwtHPMpcwI
xdTDv42TKZKvQZWhVWEc5LqnJ1wIAN3H5YrkDkNvWuyBvcEufXPuM+F0oGqvM0bE7eRPGmHpHjMa
smv4LsAxScSDN5c/ZzkI6q2illDxcJrvAE2gdss6namqve0QCwY6myb6Uq02scn35TRCUIS8XSFg
4Qvb9V1mnPE7mM1TOJoj1cMKv4Iu6YIA0BrWq/9KbHavVPFr6SV9q1I1f+fY28zPwN988/RxaBaP
pIMLIbdboUsTN8fZo9dhFgSE636VXEjGXq0h3st2B3sqkIn8wIE8JJLKK66Sm1YZkJDnRWSSCYMY
/GKSMf205wzG29a85mbIRAl2buHpBpo/cFoVHkE0FPCPMl/0TtX1q4lwvOvzXmRI7fIsGA1ScsQS
toBqZ1i/U58sCVXDL3Im2vCSMDAnVVpEM2R8ficxnQhLuHJ0zvU43Wqg2Cz3X9bQvVCLkm4svELU
AI4pbRejL9/bRfgSbK7u5pD1eYpQElB0Xx+aJmqqp2vnppkK8Ks4StGvN1x9cuoaZFoWS6n+DVZ9
m6xkc2JJ2ihce3M8VrCupadbXw7We2Fxm5kdiGIQKEac+Ict8ALjJpOD85yfzw7eCJeAIiajyRNL
K/aMJUru0I4a/yREFA3jZeIYG51TbtMzedbQoNGpm44CxH7Q45nTL5xClUAMvr+nIC5kkx9iH1yy
M6h0kJhGTQt4Dnh5KUYOQPNmJ1n1e6wL98IHqq2ey4V7MhMaOSq3uZnEmw0nrrPRCCOuadGGpOLj
2WobpADOU1NdJOcFW9bZ9FCPiFYD0gZvGfqOtXx51jpVQOYJu5LpNWfNTz2EY+Hrb/lNDpuwLtqS
s29X6IhQuhqu+H4PC5zbQD3Cc+8Zf9PrTSq2w9ze7Uiqa9/DW+Gk+RZDZIUFHLU6QDbzfvy34bYA
Be7s2VGaCu9hlE4FAXAd6AoQFyOIrw+hlGuds002qJc0SrpmPTTgf1S9NZdxTFRzJoTa2icgo0Sz
pVIpcUN1rUxzzkRwRoKK23a3jj7KXm7Na7CiBbxDi41/MQYOiMIoQai9rchtt38uOWetsmTwzHd4
NGv0h/0dVCq/qsIfusuj68CuNDCHecTo9HIj7NYkfDhTbNKpl9W9EOyTsE+xraq1kxIliet16Z8c
Iz7oy2ANU1vx6zzLeV4naeirt7WYuL2tw2OUAlwbciSl/Lu2HKOCVThv0bbhlk10lJbgY+Fp8p/+
6Mvfot6NnDvY3QITx/yKyU2QZ8GPCnlOuBuBcVutVI+3FJI+7NJD4C1ZtVwZpuodnH+zTb1iJipj
NDuFtXFv/D1JPd297WpA4cW0h3kY+udEJ9+8PvZ+QzZYILgRnoJ7uqGXsK07XOsbPCpIxaIYfLNb
07u2T+h+wh4KSJZd24SYatx0QIAI2JZnNGl9k0FHgkQr/whgxQCfiHKACTpkru8Di667KDaaMx7o
AYykc5M3TdhKC4xB1Em8hHU/KkA4MZFcigeby1pD9t+GI2ab2gZcOk986jgRKLQ0+fA1HL6+BsKH
0FRgvLq2tWFFW+ct6VwRRdsCOU/ODi1hcbl/0LKP0pyxHeITataj1g3jgB9zmJPCtbOa8i7vZo7m
RlIvc1/L3BT3yCFUqBDVbL3ZmF6mVQd2XdFxfzJBcK/FC3M9Iwh+7zFg7fhZJ5PvSqkjbCsiOKXU
ry0Wnv6uFdpz/hQA1+I0Htap4QgbUQvIWJrWFo7RJtPfr71tL49Q3nxg3ciu+iW6Mj4zQOlcrSSx
iES5b3v4tfgansRrSepV0xOWtZSWGr/0G8eR8y+0qVP1zzM73iwwO9/SlQGmb2GziZb3hLxclje8
loR6gD5aIslNKZZtv94PHtO/yDh1hb+RI/36OIaHnjA33JLXm+AwJeeBgQhsAsXl0S/2egJdD6bL
y9PH/Wx1iZHwqVZ4y+TI1QxZ+Vm7ahjDcfWLIVXgfU+enFdsAep29iDMMYPqOccuxxZ9IiJ7kKSL
yVZVKX6oktC5EpMvokyWkzD7eHAjOh/OMrY3kxz2Mfmic9lTPotM0ufHXAA/hQq1KRyEy0w7ujEs
7nPu0UKFukDe+inhOJJUHjt1xexHsUy+1zG+JPj5XKwIdEPliCO6sl5kqZhT35TfdTDKF7kc1bpt
uzir91O1ErB8OLjZqXxVi9afFxRa7GYabSmlAfm95Jczf8fl4bfNi4+Z/HK+s18ekLuBfzqbcqoz
MmjfUIq23sIqZwj1c6199+0VkAgNVxNcPeJCldjMYbZ4rQeJH+mrvTuc8TBEoJPGnSubCwyWDhe5
YBhRByEnIrJ702Y1tx1JJu+CrvqKmopJznGE/Xc1MszdfJiN+KQ+E5BhMRdUHVZsRVR28IpcIVzD
Z5QItu7gGqR9llU1LgTudGqbdzU03ydcNa50Zr+8fmjToQM24+8bcwCIZCAIoi3USN10JIY9DzOy
4y6TnVUuX6J9MVqV2sMgkP/WqS9gRupW1Cn1YygzwUM/Dn7dSCRw2y0o9cQstfVldPwQsHhcofcK
+5XDOQqLxGa9P/6RtGcvAHxxyDiDMwfyUb8CHWwLTlBAKbfS8E0Mo3b0CuFtWWxkJ3cntCnV4mjR
jVy1bUjCbRwuXgM8x4H77MqVfmZEMI5IBRs6+QasQ3rx16bmAl/MMABVFF2WP6sscgAt/Q0+7M73
UcAuE7PS7LAQ2T0SrsqDr+06daJ1ZMVli2LZTJ+Ld2p6dPdV84dvmBg9nanjSTwfo0u+6xEz6LHn
sZKuw3qh4JapvlGa32QyvjgfLNsH5hum9X0Iuk2eftxKacQu9cAm+RRhEQMt761spJSQsqejKYTq
9GiY5d4jzpyeRk2cdW5PD4QTuTaZADXZYGPpqQFNVWzvEiMvOaLggSP/7RSWIS6D1pl6mUBknhLT
8VXs9VHWbcx2o67cGrkhZNtWjRo5cPN0ZiXwMF0I0nWUdagEXGgvED8EKG82rIHbtyYu1PUKv005
IAEvuoqdGB6u8C1JzgDBL9edOcYEpjcqieu9PhSt0YqXlm8PqpTV5zeKD1a+ovLTFiHIH+p/5Hpn
EHeQKmqvuIAIs9OqAYn5LGs2qLzDfO382L4MfUSVZou/58PQPL6LG2pmFR91sW06U09oRJgp4tkI
3wELQOEKaWM5ZYVBG9ENw5eA81aCWnHTeIrHuSfGtHXoy1noLKu2QBk/uCDcYcXKTZNl1pqH4u/W
5apMYYxSvDJrpHze6ufH6bwsvc+W5CYUwaRNyeI0EGgqe2HL3V4mfXLpTVsDiTc1uuwiKLmRwb9/
F3rqxB72PUCm5FSyp7sEpIWvrjEOcy4mMH/yHI5sXjBwmNbTFurON5P9SBeL7Ywm3uoVd4bv5nPw
PftUhwDDXYP3TXfD8llX3o05JKJe0TR7IZvp7/W1HXfP+BdwbpahfvwOlvIEXI5/o5U3gCrEvxoh
XfPXqfFzJNsk7lhnne7jGKZrn6AzFbcc1Jj9F5rJchdPmqJN9LSKMuYOTcKGQPYdNaHqUGwQT2Hg
K1dfngFhTnWQEKNwpGTL04DQporKh0OMt6I0571ugM6ze7x6Kn9glZnjCMGgLbQZKudP5D2ZZMoV
4tiosJY3VO+jHYkakI8GqNQ29i4T9bYbB3SM+WzjrFlfoDsUpWWcfEur7bZ5nOhjli8NTm1lMsrZ
qagQB/yjlDFZJ4/DVSJ8vkAsqXYtGGJO0SGIacrfKId1aAtltN+paItjS9ucC6usPwR2zXn4hhMF
jAvY7dBtFeXODbGnoFjUtIG5NlodOMTcx7rLhDamKotDikSzkYPkv4XEbUti4Mu2tnTokHJ1M59R
EochTg/3OaNZNPxhODi6qEMGQRgAtWQefy6XIjNeuMJBoWtXpHaDUMGGzf2OUVdpHzWUaKqBMDs3
L79uT90k0x2evYV78iAb1BeIDRyiOiKokc+KSs/T6fqjqQgk2CrbAOIK4SzHFmvExpoxryUzp/ul
XGmvmjyWeN2xid8mURWJlLjEXp7saw6NQSww0IcUF1R7iRc7mT+7LuGJSKCfU0DAC+lyGn0zkTXZ
qFTHRQpASJrbX2ImV8s3p0EixqpmKUNfcO0MnCM64orLjmVzbXV9iaLus5/I80+tYIMtHe75zubq
17Vfi4POYPX/RuADF+rkh8RFvwIBt0l0ZrJhAPK3jrGI/EA9D+5UM1G7j+VxX0UdMhisMago/w0e
nR0Gh7BrzSc2D5bdT89TfrCjJwvtGUSdtpyDJd1tlxZHm/QqUvzj/Zh2nOOjwhFl6pl8X/ypJEra
bhH78Blc/EhRcjKIDmE35MvkA89AHropY1Ya492NGGIQv+ayS/RNYgRNVMFjmtTqWZIaothKIZq+
iaN8kDQQnrT4oYjH6eLH3ssJFTPGl1Me9L6Sq9CtVX4suQz9JlM/+sJKFzXznqEAlAXuzr3qvk9t
UKRkjONK5oSzlfzk5zs7cW+cmWmv7HqhRwER6FebBTagDBUu5j8fHlkrT3sG0w9mZpbgw5g+7vb+
otYaqyGBFcV4fb/vLGouwyiRnZYzhFX0d786MIJBK2AXgL1lHnpVL0EyDj10YK0lS31MOVBOEiI6
j1Un6fkmxttR0kbTiYdkUs1PedCG3kN85VIT7vfKFbX0dKQrkND26j857OcAbKDFMk1QX0UCOe+V
KLG/SaAl4PK0BxiFaq7VUI+MHcEwSwGm4R+Dby4DqZoq6L4qcALGp9QExrHT3+BOix2CD16+ytIo
Kl+pjjPORzIiNIBMvNwOxAuNBbfWDZfaWwBWB8SySyo7jxTgc1Mtt5SaeXvhKqXxzXCSRDh4WOxv
5gi844iWRpJ0vabf5Gzo/Tm14DKA4XR2OevNXhIHNK+EIzwJ00Sfbtx7ahnluD8v0t3q1YXTDlkr
ldVgkcPyhK6CwpChyzecVKQTpr8/+CNH96TZvvvWc8Ilo+Rk06lD95goyqIrJ3WVry/d9Dr9hrLw
NlCUUYYqrnIT6glSivXvyMVVaavWkoHG+dGdYcWHtxzbjL0HPCD3bbIUIWmzA4Ri3IRrjPWoeq65
MMDHRw7ugDwoRGye/5m1seRuOqO3L2lZNfzNvTCcBHQPyRS3qBQYILafD2xkxoUj0B5k5i3EemYf
rHiEUFVgVRCiowwI7uJWN1qj49Hlgav4D6gH7mi+YYvpBSir7I0p9NHjmbGdT25dGZ6KMlIdaEfu
+mqDMOzrdRQ/yC+8GhlDdY5bR5QbqCcXiLysDDJca9FJ2q3Jjp2+i9E6AgCHM3OBugJIRir+hFse
FPfXSK0BTmujsRKogftJu0RDFlQQlygSKdFLL7//gX2MyEwiH1TDCjKroDOrJhFNoj6rQ2VrlFqZ
JG3QKAmSDp1lupetkzntQNFwrViOwVJqft+Oq1l4APTh615s0+3l8rLYB5meLgbFem0tk4KF9jbd
VoYSgOdKfbHJg2JxNwkbhjuVzt9IlBDo5q2wYirObyN6gRu1Y8KVT0y200oftUTmeKFGHcM/Cdph
apM8yVmAgp/9buw1eGPh21HdPsnF2VT3qPQsOUMU0kfimk3NdmBEzkS6IvPaovrfOaoq4+Xx0mPA
8w0s4FJR7gGSDShIC4OP8YVFBWZDxQJVnP3RfYU2YHREarqT8YkoSMHT3+4WFCeJPldxz2mmIibv
oTlBGAKkN+vrw7rZnGlsA/ihl4botp+09Zs6CQvIzYsTAS5VS755SXZIwhN7CPzhgwHPUPmtmda9
kIdqNg5s8AoKUgq/ucd+ng0qS8OASnOOC5xDi3sUTX8LJQaQKH38WWaxoR+mAK60n+k5iJpckTjM
KdTFAiRd4UHwJaUMzecUa5HuKDU8EFJgsIxpXQYqXD3ZDs9dlLdL8fRWcEXCpIuWqlCQzbkWGRl9
WA+y6bcYxzKw4BwDt1lSJnaPu4PmL8hEA/pbAYey4GHJwQ0ZQkgXbbM27aXOT3+wGJuP7Lw9ciwn
krs0fW4D7BQ+uvIWdShU/+a6dwRrDb3vHnAVgJ5ZIczHj3V0edw95Nfvc3xXauH0ECK+tJNGWrxl
sMnmrPuQ3DwCRh/MNUiN0KjaGUCrf8PEROLZgshssolE/EhtNwM7JEOymHYkT+08j5fRuS9msl83
fAjwp6dOQZqtAe80Lx/blBOGSVfr3/7WL6b55zxgPUN5rggqc1mA2Ot+24578YxXCTVpuMaks0ZA
O7tgJpu2DfYDp6P1R1fSVboG+lQ6rDkANPNanBwhUU8h6BR7evS1uavGjFqvi9/TNyK/MeDceQ4o
4h0JAhyz6KnajWHDiNzYMXrOlh7OiOJ0qagvdxYzGgrQ+S1G74ofHBDCe6Xm2bK7a4znf8gQKhYA
8U9/Kr+YW/45ThafWrifd4UX8PvCFX+deC8GqmlweyWSTE1JRA4m6nIc1h8UvZXTYxHMHitA7X/q
7MKpqSlMv9tV/8Nv5Jwrx4oK/in+ewpSU5jpS7lKnXl9YUdwMtx9yGBNbEgZd0fZrC9Fa4v1rFx9
9wQRFPCDszMxZfxSlhPm46MYEVNKFcR3qEiSXuhDMAr950cuLT6ME4wuQzAQlzb4LOeUaGLTjONo
jMF5ZGQYjsD6ekYrdmkOs+1YVl0r4AJfUzXnZ9urhOARvj/SQREn6djESAjOn1e9K+PJseCOa0vD
rCDimV9MO2/e4Khq/YsP4X11vf8nFNU1Ifbo9XyoRsyj7PpLyAjvoByeSp9MBh1msdXVr1JMFARb
+By+B0P/moETFFftXdwmyhD1hF4HfLACgIAxpLpBOlCgENJBPrwzRjRoxSxQQ94zNUe2MeMb7X2A
RLcJX8whC1F2R6h3vQuy+5iPbcxBydT9RZ47y5Fv9b3Bw3555K+xF+RS4uYMcGS8IrMMHbzLtDZD
zmHdJz0nrG9qIM4mSTm4ZXdAOvgzjkttCrWDBW4olqrv4H3+JiyARgGYaoJ9o3LwfXQQ2NpaAPQ4
d9a72aDgZGYI7p/MKFmsFxc0B1Ndy0kclszQV9SpwaLsuSFuprNCFWVsraPqdswGRSNU3rV27PnZ
x/HHIi4cUh2tcP8TliUA6ahGNwjAzlBYmiMlx+BJNvTgk4+l/0yRKa9WY49oEvENOTiEwNij155T
15C8HE9VYU9ot5ef1h2GJ1MD+2IkrI9f4NZJ56Hr9mv7oeDSrcfui3BbEo8ZO4ynmvAophFZ8gg/
d1UlhGCSYUqFeq2ajfV2LW6nhG+m8tWuvTzLKFKFfrUySz1n53noUoeD8N8my5yv02pyp5RMB+Yv
lbSPMylMor4OnHf/w4C6O55BuP0OF7XdzM80NdHbf6cLTYwCEwtY1A7XG4KG0nP8NBijoosREPyY
Jo+CiGIn8nxKN8lTLbtsJcKWVDkpI616LTwnu22K3+gDFvK7YsQp83oX2EYfv1s56f3KerE+FJ/I
VqZL4t9nwj4iABKtSHoM3pC5cUFxVyt1hireK8vQT3DJjHWBYEXTB9sJkclPC8avsUi7ETuKZFf5
G4qIw/JR0QXjobJlO9np2/kgLwhc6haveYjuQyMVDLyaxUr+Bu6s8ZK2HFnV3oW6lb5c1hhvTasM
J2tB518iTIFICgSlzD5CVSSmFzI9Zu+L6erzfuqALxJJcR93/tJIQApaoXaQUyW+y2QM/3iBnLme
Vupx6ao4SaG3cQesjO8scOv/Ozcdn7GzTGHH2HdIOxAVpeU3MZcrPLkEAzwl32QN5v4ZHRaR02g2
XHi0XsTzfnoYQhh2h9NKMRbCcig2kgsTe6JaTHwgqI3gIz0CxHenNp7RllTR32y9Z1tZZ9kpl8AY
yCgy2Q8bPLTrPv85o0yMkMpRVt9rIPiOyuB8ueIsqFVg8hfc8kfHfayW4RVwz7UE71sUSL7vTyvI
33nby3Qoa1nRct4Pv9QqmMEtHicuO0iKJmCq2RT4zfYeILfib96Hp5ANBMA1fdvEtGGu4tpMcV0b
WX5pPyjxNWP4DIXq3zxRIH170haI7TwlT0Ua1SAspLP9/t4iaIbcoUG5ei9yVd3USnzTEfyOQp3W
LIKmGpAz//Bsrcx2mRSbAyJ8URxgzU+090dAlBD3CxsguQQ16FGtyLUsWRa0zOVW31awOZkSqrBS
y2JaR0kMdjdXruLx2NboEBWNZKYvBBPdkOkcCZOT/WOzASiiumREAUsznGpV5X8WzSf8EXtHEzzl
sjEhZx/h6zA0rlntriKZBf0pfw3iqA4N/nE+woC+dc5H4pMrT9MFgT8cK3BRs7ZzzApG1SUv0rXY
Q1FZrhdoyUK2w3lgbTZTH5XHC5SIV9sEXzKTO7Rxx/G/z0630JGFYjKXbTNaYfh5v+65S9h9LKeb
Rrih9z5KxVgUTmWdi4bR1ta6dd2t/KUjPBfMP3qDAqmjNsvnqFnKfDazmo6CdnBHsTZas+P2Gyah
MBxZXOf4luJ/a8lDtUgW3wqBgpRv80LMk4QHTE2oT6PFL+FLCdf+EWI0KOlXj9erQWR6iP1YTbss
godO0Tti0lmRlrXeJJdZOqp9JZIAhuB56v6iTuZggxeHj8hmY/N/Kb7nFducrhmG+p7lIG5+OSqg
h0arxBukfdu5ki/SKAWOLR2XVeqAM+BCCNPMHZfprbvKuRH/e8gwqA+FwK11/9LPo8LvWgah/Mbu
NYpLEMKPpJgM5JhSZq74lFRBgESYn/fGQAMGBVApWF+jvIl3tWmKwmOHtfa1AaHvssyuGvz8aJJd
4yjtQOMTYNrvQ3ChCf170a7DezvczuY9TTNZ3gN21oNT+zVOtPFF8MJ/WjZ/LvY8ExWukrkK5jLR
JDLUwywHOv384uZelMTs85f4nqRbqp3xp8NfiBbUFcghHqoFww3ChSZf5IJSwNbUgihXtkuaaaMI
EurN3xiq0zB7GxU31oTmG084b3VUs4j70lqrKfECD12G7aQIkuwGKemkCGBy64sH3KU4P81aIlyk
zpvBQytMta5a6byGeVptrBDDBGdE9rnCTp9yOH5H6pZMAn0GmtHnMTw/sEBBwSXoniW4XXJhl2Iq
1DlrNWoS+wONFp7COkoeFKZlnk7EkEFOMuZ4NsyDu87MX8nSrTZvrvpeaZZTRoZb5erXv30W5U8Q
SZSxOqwgTI0Su0xLWJPWsS9RuLoSXBiAL3+x+KJ0tNNhAaexBWUj0E/WUtGC1BlfRqexXK/BkMRk
o8XkR7JDDmx3Z0VLbKd9jb4o/X5AEj9YGjDjuU/dq8ysAgD2nZDmwQRAhb6SghUvHKCuXKEZIfVl
smTAesZzP3ozfKjYrLroJ0UwLf+XCnnxYwIpw/QiWUyhIB0fqdteEVnD4eEGP5dLDABcg5nilDXb
TkwrYMVasKc8F9cSyWFoUqUAfQDx86aYArWW8a0416ZJfnAUZfMYOvMmLCsN9UBh97ih+LBjjeUj
rMz9+Ml0IDYRS43PDzaho9JXDGU6TbnSmHIHDNEZ4hrN1y0i2nxaysjc1/DztdB8NpZveF3KsR7m
ASD8L2JBbswhtR3UAGrzz05QQ9E/BARiEzbd4wL5jAroeuWPhNGBkUckEVf0nCzYP8omROOc3cda
VE2BoDbu7PA3aYVm2jaSr3XlJzBF7RNmMvR1Pix0y4PndybiNwQwp+NVWj9oEgx/niDw626V9JkJ
qyuJnLDaaOzLY7qd2DaijM7JJrjDt0NuX4uGB18bQcojXmOVeApuPbj6EMtdezN450yzem5wp4uk
pu0m1vkiUdUEiNFb9OJX4ePbHH9A4kPH08lUsSOl2XEFBMoMNDn8kWOwlNl2fZpz0TRow6kp0aHZ
VJcawiC86j8rOsFBb5DCnXpU+rCTbsiA+HPhOVH+UGVRt70dcHbBCtV1YFBAEJFfm8ZupE0B8ou0
86rZIOGBkZoAFiIwt9bJTPWY/me6G3qMHH9xX2lFX7GJT82QYLh8ypy4WN8hC/+q5B4rz7gIVv6I
0ST1CfV6xDq2Q7gMuTEEuM08UOl4yHXwc38A6htQF1vYhGr2SrLT0ehyb1sONhhIwiZPL4jwhhql
HnUNjJyhQUz1O6P53wg3scJOw/16HPo/RW0PNScUbthj7BeSVEtnj5a2Q+QVBKS3J1f4QbhJMBv6
PsuySZR6ZosHvSYLcs/yP0a8AYvjV7tHMQfcpHPxpLt19SfTLHJNbWqywld8rrU9QJ2tZ79krM9/
I9gRuGA1eLsgIQMoKc6m9mivs56iw8vryxSxpfpKu9CK0NglDBM7KcqWW6H8IP9sjYWsQp5/mGS2
a+fjuH2V1nBx70rOHqNhjKtF2x0UW407CVDi5XntwfuXd1dQzQxKTs7UJPm8he9A9FeOMH1St8wE
K5KzhQLxomEbrN0VY1QeNTytizrqG6ML+JDKKgTcrKXGExguknFb48nkBK8+KjZVvk8Gpi06tA5T
+Ow3C1TwU8FBSGVZqQ0whN+Jv8DJDjBMPlgyj/plxTmrheQh6yeSSkbnC1KbPcEbKbPYLIrsrxze
CoV1a+F+O/+yeZtbbHpqwA5/L10MM9Naleww1T9/sF5LgWPDes3AR/vmCyMhfR0LkF2zSMmQ/Qgj
AZGaveJxx/TCKQF/YOrgQ3kQweSV/1PrBuVoFm5BqV8MM0L5WhUYJCrLz2Mssy2NhLeiPY1ORxKp
QdGZIIHp/hvFGvHUn9ZXIwcADEKoWeNPk7Dkc4TC1y7+GBI8mnNgrva0CvbEyuA29B+EBATS7ZKQ
rQ6UaPIMzENIAN/OFtFMiKdtwck3Q9nVHe6tSsRCO2ZBunvOrw+25xvmk/HEr8hS0CWPeaWltvHt
2sUtLFbzjKAxzicJ3WMBJY788idpNmXVpOQB2HYqAOECoJYZpzDVo6TNuCw6NftABfeWUAhcC1xB
8g56Pl6vW+Vha+e57J1ZpLjN2E8+fPBz3EzYrszehI21JWmodBcH0Snk6mEyE0OIZU/TDgFrRuQ/
P57CIbcJKhGrTxrvgTWwGBxMno2kMEwMI/adUAFG7h+y+t6P/XsFeUDoW5cbe0dc8x+hyPQAJsCC
vnQeX6rNNZTdtjIaJRsJCgj7qkuCazGSuYSddeQ2fcBTpMnlXnWagtnqVsNQpOgujkn3+37ss/Ny
1qWKMcSOSUESUVMvhxdkUl4toW+vhyA07CSH8IgEUjWt10suQFBrYR1pkQaZEObNssKvqDSw9+t1
rCnOG10neRnzxArUKx1uYTY++F7eZRQTlOLITlzCkoKoS99fiwwLFyt8habJ65O9AaWVU0OZKSgI
NmR6LBlowPUkRBvYlcU6xf2Btkads5oA9T2e6UiXjlzkmuU34htizTO9APk/L2a5G7+MaMaUYLhH
WVlTT/oml8Jilk80thSpnYy4xf5oAm4xal7SZnGA5+6T5G/Uy9lb/2AQEkSoXQVQBz6XQsN40KHk
jquEryg/PmZyDKBNyqOTQPQoaqdfj/M5+mZ0uNuecSd3GOteDQJQg2KPnXcEksQwlapS86VH74iB
Jwn4TZYEamru+1tfnr+bqcyIK7t7FO1F0N7yeLWnsHJ8jay4ax6del3+S8T4oAOFZuvvpYE55bMq
ileCXZOL3jPyNWBQCYgHQjJKpK0EyM5mV3ja18VipldqLchdzF7+4tDQ0dTIP9c9sq8lTgLgnbH1
kD60whXMpJoLmen/10q4u0xxnwazwfJu21yzClMnP2tgqqlmc1tLfQkBdQbbnIr6P42WxAntrMG6
KkvLWae2vpvnIX+Lu7VwWOrhpyoh4ynUSIuxBhVwGuDQ8e9qY55I06uJZz6GwjgS0lu/AFXR0xTc
TbhB+nDyXkEXXn/gjoUIh6EsnqYi1r/56idvgxLGTqWL79t6akmGh/QiRR+xJeslgINl4Y7KPo+Q
52pdyXYP3lKPFE8qE+AK23twOV1dbUGREBcGbB4WQWt2eqcpFCKol2zCkTbfP41R7gju/0uA2Z3K
WS5P7i+OpKNCLIaxVGQ+qN1izQmkSvfI4tpNfdn3gDKsASpxwYdhmSMXIeW1vFE6iZoMh3bfHIjR
9WWwlBG+AmKsQd6BDmG8TPi7MtTTNJE5dp7ZcRy8RWacieg57ppjcyyoOVkdhetZCrPqy5/Xg8SK
nZpXbtGJs4e2ZSs7HJp9QjxvsM7d6nSqyNMFKSXo7a0YT5o0RecfQDYuiRCucb5k98DZnph7b79G
sm7T+jq05bPbsfrdzwdQjmUh+8UUgJysLtRJVI5az+lcft+9kRoRGn66lOPeX3wu89OcoRIw8Jis
CZ2YdNbmjwy08dD4+7TYe/Ei+QUdGqcctc4Ar7Ha6szUCwUv+zoOlkmMz0KynmPna/0rS0Yw1P1v
1bhAVDMKCQT8GpR/Wyv5yo4Aj41YdeQm1uOPuMzC4RGsGy3lyMk29+GS7yT10X3rsxrn3EEikBL4
69y7qA0vobWssQx72kRKL/IfSIpRuGzJDFKQ2uZ+B/FxvayaaA5ZEfMh8p4ClBU2ezCUZ4L8o4MI
Z6YaTgaejprKBgJVyyHT/KUMvj5uiJiYJORX8maU8isPPGrBZ6ZYIC+rakbIXbibRXFO7+8eYopT
fdRNSdqkBno4Omq+vSC4zemDLelK2uQ20MVydSTZvQoK4HtLRA4hlaSzXRbZnyCcw27b1sMcowBw
2NEZA+vwXzbjx7lcHddx2v3PPQh7jh/hUDmoMO9fcYdf3d9/3RgDhgtv94m86O3qmJLWmooT5LbG
0LFlswzhv89tnpsTlt4zuzhCcf5SB+rpZiGW0SN5g66BD/JtrqLxPnNUW/SqU4saUafm6pqyUOGz
S6ODCNnlxPwRonZZ2AWH/ZVYoAHfoCE1MVQ3iY0hgeEFmQRO2qr7NGuUbAd1sqSy1Y4G84rL6l7Y
1/JgndNKBeAVseGuf5ukR6sAk43Zhz6ObMo34h44W/zD5jbJdX+IXKs3Z/HOBhW7kFHDwc2nHB3Q
BdzUnKpGuBFvN15v/fz63HqOaTjZYsdQ63OT29GIuLvnArC7wAfUfVHo7qGr0rcLI6T7iOsZPfs0
yGXltl0Hy+RNr2IWjXgbwAbULbzbJmNR2sUZaV1nj+GPSlQEAfNX0rd+Cw/rXIRDRg+lA4QEaI/R
l4WcbVrfuTUrn59a8h3wd809YYpA2iIfKDghADyBvWuwhO6NLeJHZhbsi+TljU8nLZS/Os36acu5
HV43ltbKCAvUJPiq3gDrwJRKZNSxkW3i5korz2eJWW6jjHE37afk2KrL2fgWWoylmDQObGF0FjPE
1uY3y2NI+ETvkWqaunEpgYjQm63zoi5Sf/LXaocC5Aso4j92w0QinUhDxUCGZvmv/tFX3iCuwG9G
nNDG8yexUMh8sx0ghoaZNo4a9v+CHqWLbXYICxMHDeBZdI/s5HICsqavB9GviKF4CcY0gkrEgLUA
GCn5M7lqqWVyIZJo2RZSysRY2G6BrTDNIv/e+WE1Kl4bohNxI4Wr3Jqxkmi4J9icKOIVJJvixFcg
o6qtrfhgKqK1oDbBvzWSGtdUIEeahyNiJDUqxT7dTzswpGhU7Q7D8YojlK/eHjI8FmyPsPap1akL
pfrggAQW7Skjcwof1prlOEmBjWgi0/1c+vx0LeQiP1lc0LxRsUkkI+vshcMkepxBVHktqUG5Vzmr
KJ48KHFzIsLVXv3ux9JNUykmlYWG7W7e9O99ealydjum71KdcPuPoFK9yoKLfgJKDAsZoOlPI49x
HTrvpt92YW9gHqNEZxe0gURwi1xhxQzX14oDvzZ532v/TuewcGGsSK03/vtyUPOAB7ZhQFbzfwqo
WQZRnkKCPINdz+3RsDtY9jEfNpIxrDHrbA5Yy2MZEW1dfFtTBrp3NH2Vcot69J2EXM149Ur2URzb
l4DZzm7peZwKQnTIXmN2I19SN/exaTDs7NcE6PvHEDQU5i1PXBTopAe2j+wQOzuGgGG4/TwO2JLc
92vtKeG1WunlPngeFyeNwiQjToYWj9kSKcyZsqy+JrT/5rNVb06irH5e70EL2j+It0doBTPcF/NC
QSG4n5qtZ1NCib79KEn0j3mf8oJUiLBx6wOFDGHdZiKi25SWpTYM3MobbEmG2hhqk8vp2KHCwSs4
XbSszsB0VWfwFkGlHeLx2Z9Vf4+3g0pPehgpvOzY6pDgEJk5zuPYGu6PLkv6tfNfrbVwAf36RIBr
Ah3txsZNkZn/PLnX+2wnVlpIvxMcYCja9f3giVDo1CNlv/kV2vTzHXjv94nS6MV3DdhpwZ5IPoB3
Kw/KgplaalpuZTpuZnCSfK7BZbN8yeaZIqGfRbLb7ZLww1kxMhl8fzIaf9WB9Cd6buo6ojm7IxSf
Mjlkfq7hulRJLeHrlWCJwThxG1Q9URuS4mm4W/mPyS8vY48IZ6lAlHIfFE0qPee4B67z/mC+Axne
QJTsXpzHqE2oOrREI8l584PUxoo5nCIdFjaOkFXyt+x4yicqRZKrfPUlzWCUtpF2+fdwFtmMdHFW
rVpf2vugKHv/n2H4Pp80wxm2OWc0X2V4e4Tau26d+qFZ1CRs49wQzQ43V1BgqCawe5YbuQnajQ5+
m2zN8LOHJOrUVRdbil8B3ntW6l5i/BlUymmK/JFUp4m7Zm5SVSLHbya7ZwSEz5XOE6gchQD+372t
t/5t5se0C9mAnFmWeL1XCnN9Ko2Gzb0Fbim4JIFEuPOQeACk1WdXH8jNb2WsHX7aPYl2G25Z52So
KP3FKfoBC64aJAHDwbTFT71+97o4xUIoN84riRueET8c5Y5z9OigIM2yxf4hwDTH7sfC0UkRsztd
+6SO+pfDv331vowk6SSFOw4eh0k1ecoFyjFmndmcaTyOjNYpGyj/RHwVBJVJz/DZaqqpH1nVu+i0
nQ+NxNQWocF+gxcQiX07m2eUfVO3fpVRP8U9/hgxNA5woyGZbCmzZQ1YjED3HrZD7X+RM4OpGtDE
FKI5KZvy5m6WQ/XoX8PexedX8NmRVjZyz5swdb0tisiY2yRSeJDos0N7CpLtsgkrEx5jUceGTI0N
igIvDBrqqDMDCaVoW4CLcXiu3aQyPC2evJZWD1K+NRQjivcjlmq/hRq9y+FIdOr/MgifPX68SjFC
7OfCqzyU4eXe3rDYE+aenTpi4yh9T7NOjmhb1PW08p+zozHlnoi2RGGOTUdalm5kP5Cm01xxgNhE
X1hvDVInv2xsDj92UrDa+HVaUXipteQ9+Nr/L/+xxpAegjk+f53gtAu7cnMqs5hOu8SCsA/q6R2g
Re9Yqh6DTRy8CHiVHboDP3NEU9XOvnXC6GYlKrZ8PCFm6KvEC5qPsP+JL99nywMJdCQaxGePIhTt
ntMyGXwp1DOakIXOHPnzVo4cJ1MXHs3dmHOe5qOBsLMswiTR6q+UwCI5UbFT4JAJCORUsZUnqeMQ
n1kknww7fH9nplKJxvX/uN8cQPsyDoeJztsapROHKlIfMGdArp4cpQr7F2pw5sIp019Cf+bx6BOZ
PQhc3nH4VlcYQZMcJlbtiRi7H5yaIQsglMsqPvLPhozGB1u4WcbuDVi9N+NQLCg07Sf966z+ASyU
/tkQdhDuhBxCJ53jgL2qQEbjR56DOPKQXNkeEZEzomZOGmifYbCkni01jtf2STqty++G9P0rY0O6
EhjxmqpJrQ6dwFF2UyRczgwp1WRT6oshWOOx4n9JMZOC4V9+x1LvECD3+ZuNccdzHDrfbsqM2D9a
1VqV8BT0DTxmqShnWFhUPcsqzxeDeH3pahcwWIrYXmzE8V+ws7APX84H/NuklG9asqxWQq5kg1NR
r/uTF1IO7iO6dvCER7aoSCXQVdNIT3KpkIcGZBocIEXoDSXcSTXi99JbIVSquTTjFQQOnQvgPsiC
1qQQMDZzh9TKc/b9uOn8lyAkvIxxTdZm62cDMNaFzfmAzOb9ZvIc7+dYbErrNO4Ksc17kq+TUW4J
+JbarTmUAI+0z0wBe2DCs/xidlMNedNxPoeUH3HSeBcmdKo/PihSZnpQreukfRKeG9nS2W15/5as
bs0g/ZAmG7G8ggUH6l/IWWr7mTFWYCRew2YrxSqok4Mp7WKlA007Sg4XD5CeCVjpWkPIDqHrOzEB
v50yUnXWTuXHPoret/BTNib90o/RprCF/tOeZXPxLgC9prBbjTmDtprLeDwxoriAC8mg49sHwDWg
WjBHH+CZGSMjzV18vrvzX8CBxQEh4IfaaVGDJd2nfQuH5HVLD4eEUUASQ8R8GnEO36/cxPLEopBg
7r/gzusRcmd/VQQ+xTyAJ1bKnmktiEpxfKypRxFZoB/dViK38xH8CBiRSrjDsLNk31PtDQDzlXeO
bV/svl/aBao1lGQddZn4U8Nn1i4MGkqcpeP6B5YP939xyRevS5vPGp4ZzXWvWBst9Wo82x6r5bRx
xF5lKc8P0/5fBbMAA0/6Wz9n7h2y535Ud3Y36wjDR6G3u85zHmvm2xCJbOVj1Rtd8hsi5E8455K6
6sLNVohrLl9mpChrgqzwlq2qhI2OQaBHeL66paTyQ2Y2sZ9KExCtQmnm3L5fKAuz0i3gHEGg4Gml
q5auCv36/GDeofUNHISMyHyX/NbGeIef2yQV34AfuuQt6fzrNA5GK2Qya55q1VSNK3TA09dntAEF
D3qe6HL7gLuLm0ZQ8449duM7sLDNSoOwWw81dQlEVacd+pKSlIJxJaTUn/YGpDuBXqEwRkuHi+p3
zsUVkeQxrZWxlInuYbNKxZgYRVaiidNQbja+nJu7mBKIpBP8n6yO/YwzhCkOk+wYDYI9M05Zquge
tmlQKqbYLMx1XHIDPLfBs2Gl2oYfydgncblPAHcMjZk6t9UEJSROkdMLaXHLAYCR1bn5mCYnkRbt
PhOFgkOAt+08ygRtuwoPQI4u/0CL7rJqq2yL0qciMiBDHyb7GJlWZrVDcdKXtTxq19hRomsFA0lu
rOiYP9QQsGyPE2iDfP8mYsz/2AIEaRJ5oV19b3nCIZdfod889x7bqHqShlbzA2CHeZvCXRWovxcw
SjPeXjfe0H3kA5ZA+nEi3Bc0k6041lV3JjB8e2A/+LKjVHtIq65Djx8mJzCYZ2KZ1ZezLk1VYFA9
4r/qYnzSanLL9pdlt7xcXludmc9PwwYqao3ifVPsV4tWrxEhugg6iD2Dw/FUZSz06aPGH4rEj1xO
s9/r7isFfBvSgMSmbQq/fx+H0xmwHvknyeJRGCB8NUo3Bl0IAAyASdwsRCsTeiWvh0i26FXi7yX5
/RscuwYhqXatMAj9TY+mlfWUkPKlyaXj4c+pjLbf0FfbDjrLH/S72Ri9SRKC9a0Kubs47CyFWu8D
v37UqP94cLj/fR15mADonL1s8GZrPu+b49Tp6Ez2as1Yb8+PFMT68cxq+BvRm8d8TlbEZX/AiH9Z
oMF/P9+SWqGNxUkyVVG4aOl0wC+VUEkR6w0MG9mIykHWC4qLm8rqXNjCRJ/lIHPWeWyZac4U2n60
09E+wjeNkV/mgGAZWo/RklQadn8lZ4OQr5qur4L5jnhEB6ZltdmGVZscxVQntWxFHaHe9M8J7vPQ
z1Kc109KVE3eGSdi/mmusq1DgsAXo/MMsCZu4fdHd6S6+Y3ZeOg+M6UlBQHR9rt18HhfCFq0MnWl
re1LT+dayFXn+ZZhko1mYybEMNERWggjvGFLe59DJgDAxEzwbQBghONYgPNIEAkdvQmdqNtQ7rIz
I/1m/Msjg3oRkPcl1yR8VS2/96heZs8aMkfuI8Ft3xkcM80RBveowTxKihJQW8G3JVX8CnmHijwl
dHzKbXt6ngJWkWPVK44A/fy06wpXRuizS5j3Ja3paNmdqXWkopFq594sd31MzXhTmQh/4xV4oAnp
Y6OPFtJIFPKPlt7E5Gm7BRsJxU3jvAhzMGkFv/x97Y55Dg3ujSkP5svqSi/SlyI2qkr9OYt/jk2N
wuhn0zHpg/JOr3CQtTc3cAAcmwuDbVIyfk0ZlYFrvY1JkRDaj526eVcqSP+C7cBJ+yDEyz7I1lZ3
23fM042hIG8LXkd6LvdLkZ0Pww3D3bylQ58ThxPA5TFevFzY6eaRBp+Z4+dMipuQ0hqEAdDSbRFA
QjwoL00E29ZxBnd3rk3lOfyFXQUDJos6v0DRUOWApbWbykyXVes4go7FF67SZ+eN3r8vocTVFvFP
jzk6MZBnLh67NlqsfGgf16LzZxHJnHQ0NvSEy2yjLEEwO4lyvMHiMPWx3krB1GtfntejCYcei9t4
E8Pzw0SNyJFMtKJR6gwWPNaRrti94id2Q+Np+UuGetjiaeTrf1BS5PgZBYndk7e4FtQwIqhpjR8t
l01Uyv1uZpK3v8cGiN9IFPHe2K/5P52Sqb6vayCZxzxrO6sa8bb89TKICQu/Ebc3aiq+tnq/A0nD
eC+XQGF6k7/AeSRv937DoHwuFYKqNIUv8ysxcEjtaJ3NngjBwSB1ewNx+FcwMuMCYjzuogvPlACX
tIy24dfVZLzd/4DGyi20WMShi0SJ4+iBFnNuBw+9eB4Dr40D6L8XGjc7OgvtgQmBzXAmZfnWJBj2
1tDNT3AWMnoi+8BsFFqAbRi7uUskfHLmpmYBIp6bjPnEwMoJEpN2N7dFH+1l62XKlZGW305wluVZ
glr83dV4pOnyJNx4IfOmSWQz3HbVBD6X1LxdVuD+/dKTKsSWFluw+tzHBArJcwIvLyrLb0B/omsN
EQLlif4mbI2tZ3ZUIOwMA3EpkbeAxmROy+RrX2DJIuQycPrxQ6Z8OISY419u97V3Z37Wl5IZE214
RM4GexEYyzmB6TQDV3hLsUUSYrqXUn9T0YpMlwx5Qltb1Qer6PxlbIJ7o+jXC4oeJGHuzXJ7tF/u
dYHs8X+BM0kEpdd4XTfNEyIeIwFQUEqmO006T8orIGuj5y+n8RogKOrVsTaGMPR1gSM1REmWoH6b
goOoR8qHeO6OCAW9yw8rZEJ57aDGO6+mt3iJvQuwBeak+EqR8V0Gx5j0ZOLexJg1/Cr8htx/iEsi
Ia2xJ2V5xZi+XPwc6dJ124wqNGJeNSi5Jrd/yAb0L4flHUNeZZaqMkKwLhBgUjWc+GiCElihWmwX
QOzb2AIrTyNJLvHNObWwDxQUIE8dc8K4ctEzDMCInLKTbK1TRlxaYVuIKi35siLY9egAK1L5ALrj
q5l3pqqIPt3nF9L16QWeF4ZtvcuSm0mGcCrquRCFndCp5Gspd/Gx3OBLf0Pfhi5FZYy+PGi2lImk
lo1T57sqzG6Gq8/gsPhy8BvtKV6NWVnqxtJGeH5SRd/uKEuMP5AuGpkHic/NwzSQYSiG5ZP3iETR
1sPFFhQFFCOzRgW5Ksy7SdeioEMjqBpiEa0e72YkfVJ5ukUtbA888ZHMiPxl6g1gLlczfi6AegDq
xS0O0FrqCWhhbkI7kPHK5st0FWemlnWmz4UieaexCc4c93UZUp3Sw4am0JdaVr3XczgW/sV8HTxn
en8syjkbmlXIWLZ8WaxTfQC4vjurpPHGIKX4tY7wS8J7pLl/9awEjnsIREafFm0DbPchr4bn/sX4
/oDBU5qwRHh6BvMkSGlGHkI5T16Vq42+FW9Y9vqHJJb4h3GDcaWBugkOaEEYOsCXsEDko6thSsWi
NJUECoVvKnAkxEJUjS1Mr9+Zf95RcYWDlIK5MvXIMaJOz9IiqWR+9nipMeRrbh5cAcvFSimNU7mM
S6dQNEeGjmrnkoXTqtObMsNVaonGA3aT2B5t9AQr6wmWMIq0d2zAokklpc8Asg17FKAl/bzzHfZT
cpqJ7anaae3fbRr3cgo1g2ltLxaAZP6bfNWUlzoi2JCqNlXZlVPNhjTvBoPqYtgvHz9UC+hOe1tk
smVEMYA6RN9pT+0jHryBweHn4ZSB/lk0ngCJwj9mqpiVaSiDlT2MCkvMHheiR4+jVy9zRVkMlJjc
4M9yf0/5pIg7zhh+sKFynU9bomLrOiaX9RzaJrDVLKvEfSA1QdkuDEYP3Gw6Wph3e3As0LwYQ52e
5HyWHu7CRVTlrIQBE7YkxXMVcQZFaJiwdpNQ2VLb9qOdRLUbbCfbac9ZbcyVclLvpWDG8ZE00G32
858HYx4SNbaLjUNTBkUVl4UqMaAFBNMGT4mf3Kxo+um+iwjnV5kDvYp/pw279mNFGBht1FFL7iVu
t0uF8xpewGbV6IYL8QIgjG//XGK8tMcuw3f+id/DnoYz4oQR+qYNiiculnsREwnmA7aoyarVR8bU
h2CWCYM0zK/Kqg+px59JBwwFN6liGRfUdD82W1LsPfxxaRPhfI2/3xMCFMg2EYkEPNshYIJoHa8w
UxQPJG7U73YKLwY2AuSh0Fwg2eJVIeKQAfWD0CgQ2vhazNppi7LDFgZprW/TUFbSlKsjX3WbINwi
SL+KiApCqAWAMYMy9jrmzszl/HTO2wqQD0zPrq/iwIRft0BkFh78O08y5I3YFJ2NsDDg2T+2OsNs
Uqfxswnp82hXAdkGXiAoTI17/f4T1ka+Qu5pHcpI6Yn57U4sWTPoF503w0W8C8xoDXxfjjln8DJK
oi6OfzbLnrMf2x0YR58MOPU7edvzcsUk8WIv6iVlF5xTpV4FD4Ky4NQumNVEi6dbV7IJVmiuJ1PA
DFlrCcXF0mVUCFv5A4Rr7KnViAtDmu+kXbL+/Rb9YdggcGQtm31Oa6BONeeqix646okAik/wY7tt
9+6SMloUXeU24Ft6XLWNQkARH1eqU8p7iaXRhRIx9WMr7bH3c4tZRtYyLHY+lXhNSUDsZKwXl5yZ
mwyVAeJyZOtX7bPL65W59z2Svt9CC1keQ35ZzwbM7vYS9YHIk8M+U1Prd/9lidzLfiA6GVsHhDLG
NENrXpQySWky283DYfD5K9nOHitJuFZqCc71tT7kkfJZ+Vh68dfxclZK3Nn+hyiRsuwAX2tmur77
cF8YsTDNGty53YAEEQcofelTdSoEVAaW5hxsfGv7nt48RRRdbS3SRg68m5d4fHBo6VvIRtMcHHvS
nl3UWoqpYiMNzmCibA0ovuZti9mZ2sdTBLZK0IMVEHM3Ws/mTgfxxzMVljvIj7kO6a77v98xQiF0
vkOaHmgrdQXKM6wV7pQTa0VROm8VditoEOkZOtJsG2GovY3o6H/S8aJG3uIzUAerG97yjsy3rt/8
3yubmrCqLT+G9gygUg/IWTIpbziKuwvZMQ34rr0glZmCLbMpcaUX0CWMEp/DOqJVCYawkGBLr/So
KSHmcqfgMtHZiijokk9F+WyN9d1gCROhRQ1fiwE+5CGdATBRRNQ9uSRJPWF+ki0nIo4N0icqn+oU
qLLflV8G8/wtDKtlpFP+8avq4GK9zwEYLdW/E8+zUtyXZKVUn4utOIMoQ5ihgvrV51eTeTxZuOvF
XpPJwycNAYRM+XJsX+77m7ruLY4m4IuMiDWk10yxMSP29QuBRTU4RMT0tq39BVwIe8/ras0Vr2a5
+lZ/beWPqO39W6qcKg/3N4v6hSiMda09TrjFxX1C63zfucNh6gshkxIjMb89TeH7nNLOs62WobaF
+JSxH3nv0YwhwCYBO0zkl1l81RWfdoB+upm2DbNmYyVPqXLopROr6ds3cX1FAC2Ntllo/y0tEqZB
/aPGKaDgKHVosHWb+YyrQxznU0W0xTdBvHRrQLhjxFoss4b3CX1ooI+WMcFGFPT2CTYWIX/dk96T
0bQGB7WHmH0WlBwryt6s9gbxxtSUddN0jYDvAiyYd3i3RD4kX+9AG7vyuQA4rEJob9KTYKDYT0/O
jgyP3YXT2eTwzUIDmLiJ+X/qZkxg8qdzTwSg0Vnd8q70crPY1zr64uo6KQr+FS+rMD2jXKconpeB
BzkGx1Q9xz2sdKv7i//La0GPc7Hwf+13PW0Mb1f8l6CF3KxiO3uM2anZyMFXW9hlvgQEHluOCu9H
cjeY49RebDgIjQh/YHJ8YegBg1RXVFd4RnmLFhJykGTr53YZ+CeaQZlPVSKlMt3SnRbC6vCROdbc
jwqJvUPu7n7BfhjZJNMKgtC8eJQABxk4EmwjpWLOrbemNYZpftJPSvXXsoy8eRNfj+1iHkE52D0L
6IuIuFnvJnXy/xJ/5qChGBjFT/GdN70yNAszHWxaHoGe8ZLHmq0xim2q9MGhegOfwXJB8O0p6Plj
5SZ/hq6TIXywLfcOkj4VtQDT5F1Ucd4axXSWB00QtNgrVvVojqxhH437DN1vOmw/on5KbGkJpta5
6eaXEQ6ldsHQBTlWYKvXg+MWH/Dq5Fo6EvMGzd2KFsJi25TwYSQ2OvyqE1UsHXMaM9HBy2cyfyhx
BdnlbUWqev+8JkhpdDD2lzxTYP9kd1VnomHngR2DnpAfRGQwQqHB2dgUUE0yT3UNGCKHflYL1K1f
VPKf8hBXkni+VtPpbNtlI5is2twjdn4sXgqeC+OevAtHEGTfp3o4RlvU3K5XqGToj6S08kZMUwow
/0UVZPAQzy5LeFUlFk8er6q+KQPQwpb+wWfhx3P65bV4XowxGF5FYln/sfrqyY5pm6gppO27B/SO
z5BgUFeZ09b7HoHh+vekRX15RcGWnReHd00JZcGIOrxJhmuyPhQigU+i/Rmvp2pCgu9l7mEY31TY
l6qjbsoI6u9MayKYLdIbOJ1pSBd9rMX3cutDOMOJO3NebpmJ+8j4zr1EQGAv2bmFbxSWtRbHNa+r
MHcH1CCORtw2E/i5wXlDFb1Gfp4OjnUAm/CNxhVT6h3lzJ7wmNpSS78UtuMvwlkLqvG+wSiTDELN
XXKzdf3HvseMltOJcBs2aHHiKjbye4FIi+gLnijgW9O4JPf8SKBlbvCuYd2+IV1YazCj7JsPCDeV
k46jx3jaROQxYjNMAlezaDRt95FH6JkiP2KFDAsdCsoD4CnanzqGp7n+rXiah73BrZSagmxbNvtd
3sA6UVHHGMdW8Oiys5UeHCmnxv4pbpisEb6pFkG7rxgWfnU7wGdA3kqnGUwwM7jQKCqSZwOwXrYa
+7VL6KwbVRh+TZR/B1o/GdFhax2Oz2B37RuSGG/7rY3gApiiwkf5LGKyuEIhpwZG7xhB+V5yvlCP
aW/jx2sTA/kYYHMU/WjPFwS740O+TxnVQ3Lt2g8KsGLlNA8nyuM9xT598am+qLceEoXpsBJDOwvk
ekwFsWgHin4PrcnJgjEhqDiNzlda6+5SVHjzdRJRCh1dCzBhoWzbTxABvCVKsdci/W41uvsm1rNm
3OIO58bUGi1FcvfABRjE6AdGT2a9MNA/MO5ewClLhPmXO0MENfc6m8u658EJfsaNlBZ49dW0rqSd
bcNARQBlwTh9xrOhsVpuq13VDEVk7WPKlVgmKILmrZ4DLirJZ1QdZbl/Xa48ZwrFIv1fvvvaLDkX
m49ymGg+25CmkYjrlM62DE3xqz2Mn5/na+zmyo17304I6Guxt0VJqseTxxNmGbqdf/Kw5GiYdZUO
YMDpcP0qLrrIDYpqFe3xIaOBo6Wu0r0sff+G6Vu044lBIPcMrxRhc2bR1ziYE3E3lJmVgsQuK208
7Iy1RgpyJaMoW7aTHkP0J9qIDM4UzfNsnKEhxujjYhno26W7drlOiU5cJbcwOL7FCWpwq0IlkkKC
3NW6yS5zVfzVJKide4VmCnqj5ZwybOVpgUUKD2VTje1Bx2jGPeSH7FYg4crqSs/AQsSrj5OUUE+8
wVztGJMH7NGDu120ozVt9bTIzeMvw8Gxz8k74gEHs+XucSvvw8vudVQBYTaNZEL+Xhy4FZOfyKOL
LHONOovDpmRvHz/h0iIMudHruNShTPajkSc4b1hvyaQMzeDlKr/Eaujj/iV3aLpF5FC860Ckujw2
0s1pfqjvaqpV6gZj3i9knQrz/BfwwHnRUGHixoWZXG2lhWrG35DijT87x5fqLefUatig7E7WTie6
ZRHfdtZesEqkzE6XfpLt3XCsjQPP7ltLd/C+I/8rCBD3wfyYHOnToIeE4MdfAXxZnth6YMq/C7uG
8fcRf87lCVAKVswZUh6LGvOAxi86yBlnmr4YiyomDQ7xMhV8NZj00NDcwCsfnGLqScXbl94paYVv
2tgyGbZQHltFvsfe5bXQp2/BjmLxdcMeUG8NsKqhW8dV3RFOn5tvc0D/3QBd5ZCAU2bdRckYTEBW
gZjj9vXZ8kk3GBQOw1SIYmvZhaabCJ3KtXvSEUVNDRlur3RVDfRkvjgYhgBihuA3bBHRL3FAKvoz
XYn2wYh5qVcv7z2eexxZiY4sMfcKBBXJ+yV07v7JtOH6qKMXgLJXf+RNNClk+YfFUw34bear+5Cl
ewFXi7mR3OsBhsoT64qHWikbJdVHG5JvkrHZ0NXRQSCh/RrI9r06KrSPswD4yRR/uy7Q9la2iEBF
swDmw8KzjspUTIxZkleNrI1rNrlqihEAFnq0utJPUV27uC8rxrz3hQqdebga26iMvWHu/UiULVvN
MTwNy3+eWHHyFVAePli7QMXCv+rF9sPE4da7i1WSKDwS65HUNCn55bJP1pYVXrIRiX9ONZvauU4P
rXjv7C6XzGJ22m7jJpp/RSYrrfa7ewUfnR6brdL16ps7/0JRh330E/RloaYAV4m80L5QTnHpB5CS
kT948unN3ALWYqiZRfJwRixE3WcwrZSsQokIJXRaxg+/pHpjG8K01lYutHGT10OTjpwihEVVIIn+
SB0YiFJQF0RCzZzy7zwhCIPB3gmyeXl1+y5cgw4zC2JYKPtktqIVSSXyRY93giyuE54NQm2XxhWR
mIRHdsz/5COChKc5fznwFz4XhAU5DgcvBk/ywVOQrmBuTHltkf0YBLeqb0wcyrdcgZ/59DdPHORX
7fwOkq+yjjpjbzBXnkYodIMENUy/7rjU5jf0gUy5RFGRIpO24Hi5TySqEfhRP0AxPdHAiV30ZyKA
d7/sSndYMUuOGKdv2pN0oUWoeM5xL2lqemsawP+RXVkDEjz8hnZde9RQ/icde03CcaEp6hnBFTcP
496e5Onl6MCKbGwwuDPyOXJgpVoPbckGKQ7rfAXmSQpKiYdhc43GQS/5IlPYl06vnI6FfLJaYSSA
WOsdBdKPSIE5tnzFDMt7mqWq5/Gs9Ll9nNAZr4qwro5H11nhgpjOzuLFRFLXX9vzpqk0eCYZRD2b
AqT/cGKdgH5QrDqQDCv8EmD1do/5PQ7kNt5mxaIhIdujJDOzhOm0UeAxBhIC3MtTS3oJZHO9xaU0
Bdxqmy+hbqOnAxeAYO/M8JqzItIkql9P/TrazJfOgzAmMsx93QS0VSvrxvGyHz1bSM2doKTxKFBu
REdikLTdDaXahDlLu6Ht4nl53cGMa4YKwtaBfgirpE4/cLRBVxJ8R5kqDGRa+oozr48Eg+5pkMqa
jsr+D9ilL5Fj/IcLxN8TRm7N7Eb2It2+FD2IjfUkzNVtGmwYbKpN5/OWFLgwlyeClCdSCvX4miox
877qDM/5w88FRhcl97Ce/mGngNG8GYVDHuKjE+1sKcyzs1a2ert5sbOZ66N3LjtYgiUvIHIIWvCq
/SO0VQun69cw/t+fGjk5Mmw9Q542Ew4o9oFRm9VXnw1cCTqnbvbe3U7r4h6cTFw9yWi9qSRULAku
hp6TzRz7Ca6OTZMSi9I1ZJz28+lcjwthRcKIfsiwFkcVjRa9xdwbYElJph/jwX0Ll1BIZ9mBvU2u
j9rDCS98KepLVFxBVfLfqKT9iTABrSzjNMaPA22TwWb7PTYX7KOWb1zVgfjTE9oApl4McLkzbW0P
0JRsmBc+BQmJf5pB6EWqpNnXSi/5Vxl11jHocShOvJMf6HnP84dwBZmAHFxqjW0gHKqaVgYaDPXF
VRqX6KYEyRu6xBBlRSJJ2s3cMhdeDQir5oXJ+K2eVT9seETiyAM4IOC3hNsI7lX1t+syscTtJhRN
5xaJdyCYOA0WBsZMdOKGiTDFbbXwuLIXuKGp1c4oI9yb47h2alrYLJnc6MgHOhwdc7jCPutw1fI9
LEpbc1eg4iAl2rLslDScTefF01YGKYkfZf4a3inO2gTNpDig2KrWBeUxK1F/VbXAcnVeQqR8axwx
Nd1PZzfTyD3XGIAXTojYA+3e3D8ZXmZPj1kSC1xLZJqkQcCUie+MwDgi9F8XaK+siYvdaAP2JSHl
UByFwI7CS145s1Ym3pTbLi+k+buJNAXX15xgHnYU4m9gWNIb8zmaxUt9px2WFzuQxqPDJa1RtJR0
zjzRYSklNIoUj7YW4SHe37dqA/uHO6mjJpO/xH1oM1cYe5Hh8RXhBBEiEz24lAiIDjS47l2TRQMy
bQ/A9URzfs6Z21NMA6CzTUV4RRJ0FW6dmWJh+4dhpWQjJTzPuBDdhSjDDxraluFDsy8jru+0ikeJ
A8I3caq9uBqSsAUbWmrOBUtrN4SEQuytJ0OzAOzJhkOl2z23gSCj28XggSKpHHGeNEfBPZDtZyJx
ysj2b/5CykwYHMVYdT6oWnj/nJiAoHBDLbML5NFmpGI5AeXP5kXNk1mpCDdhEuZcrQrwl0SZR0iK
VczdXhaLURYhPZbHHVaGWWRQ91CYZA2Y7n/sGi7BQ2EBmshO/nHezCJZMUcza93uT3UjofcmE7fJ
13veuiSRut7DpwrbtSHSNM62ltykBZG3vBVM9ulACp8JH6Wifv4SgIIy9cuAkfhACArkAtgXzPx6
hL+sH4VGG7WCOWIu/LjCTkEw3HRb7YEsj62DuGV4rVMjohKbVxD3O81NKTQr72WcRqXgJuXGQA+l
4g3awNex++LkRx1zgSQGPs+fBMlTBm54K6tneiA4rl/Ujoeb7qUgY+e8Ut8UvGHKzRum8Hg58/Ap
nRKcimPk9zl900muBAXMogk8+0VpTBKqQB/sDsL3OnsgvpAxBwH3POYN5yStDm0ipHPm1bNUPRDZ
pbn3eP/ub3U8ddeW7aFyrLLrcKxKUtFUo+lnUOOJDGrp/kpZBggFfp/PAl2qu1N1rTM6Lgc195dx
d7AhXPDNfrSqFaFXIz5Y1pB6GQMkeSU8zlM/WJtrxoVKlbgzhdqSJct7FHJRHV5ZUMf1KxD37aXA
5ueQacubJ9cgavmQQGMLHngpYAwEDkmfqadAic1KHsG6/qgNn8FnKXcrmvywALcRJatfxZH5Prfe
735cRIL1FGvrdWOp45uwOBbi1+Oi6JkNEvSvdXEVtEfcRGIPNl5+fNsXFdLMN8XaQZ0m5V5uc86c
U0AjDR9CC376ec4nPQyeeP4eCuHgmrAmZZmzEHS5rWLkmmC/U5SIvsTQ5sW+Xt7p7zy4+ISb9KVG
59ctkjDJg/qNDQ9uHCOQd5nbJk1wmeiuGyfxQ6t8TjBAaKwrNAto7xcAzx3ZTTLsiWFPpZU2Nej0
2JfB0DXeMYKWZKWsGzJT+fwEuQXkmsdx7CRjXCu4aAnKlMF2SERXp9EBXNGuU1qkmUGL7kxTDVcf
jKNNVioJnjHawItbC2ZO1bNjmSXlDBtGuU1eejGuVg5NSNbTCu8IltS2aKV/gsre+T1GPahBtRHF
WgAa8W+2PEUhSUnTbzenwpTqVJYHFc2aYWciQXskcfdt/W46dBp7LiaPoSJ91SqRUQKjeoyEc+Sn
s/x7W/UwI6sr+YDM2tT6n0gmqSpl/MWlmLHaYy/ejLukM9XW1j4Oghw/s1cBTP1BsatC7GV+1XHz
pSkDUWSItM7+FdCT1jK7fjO4uYJHuZrahJiAN4U+F2izfAm7M4+9EbkZS064h+WM2wRStVtd1mo/
9tlF1tRCdKnWEzetaDWaRDDmPkP+CkRYrc2J0kWmRdjF8JS0PdtXsML35iSadSIcZCT/hFW4kIKs
fCyW2xHbS7szNIq5ze45Rke6Q//+VA9974/JO6QoTDa7wrNHK12+ejYv1JOfeMQrtSsBY3ILlLuU
WZ7BOWPlaTbMEODNRzdm/DwV3jZGG8Spx16vIGzrnof/sAcGq8s9duW1/91ogQ7bVRzEIW6+IjKb
JvZtbY/F2bD3P6geNhNqBfIyfzFtLLVp9+XamodcdJYoo/w1BtgB39zyDpkX9hbeGHRJVRDKQAuG
LNoGScKT5pIePH7brs+4BncrnUInPh/GQznAbqyBufcfYrjp9cee/lf+Xryavk3bzCMy93Eysni1
jD0LKgvEgbZFfxmdl/5D0eaXMHd9idwLp8JPDk4Q7kwWSqwvbxji45vycZaRiiHJF22fqskKwPlG
F6fGFrUmlZHGKUgRDXMvhckkmGGlrjxh0s6MffF1YVHt/YJM385mf+7OgXWPBNxCNQHK9a6kw7ds
h+wUaRL6WaAgKaAOWGR5KEvThZwmOSDrC6Wg9q9RkoZXJHJTjxp90PXiZE/AsrBDmqqzKP6qEfTr
bRU6wpWu0PDvPhYTHCgCwdDR+/kIJF6LRBsd/p/qGTgMg25Ja/+slqKkfglWuzBjYURp/EJ/DGEC
Wkm3G1pRbKaqu0RbY6W5qOKT1uBdIkLQ88yt+0XH1cetnfEeU7ILxoTPtGo3k+wNi15oCaRD962/
z8lo5w3D09vFm8SJpDXZ/GinvxIpc4yO5SbPKF+m3lYQ0X6y3qtmqyjsSMo3+JsHlxkjRn8UTMkE
bKXnySodA6Fq2Tz29/z0G/tNHHQ419L+yIem5DHzLXy2CZhTzgxowKka2RCnk8+VJ2RPO9f7LjMg
tcK7H0dFZfkhB9o4/zT9Y1FkKpix3van0jTuVBKhT7ub7yHV81T2OLgL5a1KT5x0L3T4/8nnY5ji
69FSF5RkRiEEQZeM5TK9aLtIK9Nfis2zHjDm0I7VTjlOqtCB7usJffm40VtBJj4XCx6RtmoBLwkZ
qdSL8cqawScX5khJTfKDKLz3d9Pheq67vsB0FMrGy16/+cbeACQdd12FD7qkELAA59h+ssCabg6z
DgQWBXHuD/g4MjxC0Sysi8mJvcg+qLPWJDKh/RMAPFrgJq1HmZvxUwkAhUBrZYRzbrVoBp9Yt7GJ
VmXZEF3VYoN8QZnLdlQfTiCVegAM49IUVoJ8WfT4tR/S+NlQ6GtU3a2cOV/cJ2ZXbI/5es+xTDMy
/TpJoJ35oYCkI2TQg4FGve5izj9JYMJvcnZ1F5qEqwbRgJnugu4nraMP42dkEoN0y8SUOIfCv1rv
+iZbHBi5cUfVEzc8hP47mGtrm/jJrh9jskpZbGi6y+g+2VjPKZtK+Z75CpU9MeJXxMdSQMZ8cDn9
fCWqrEdCzdNy/yFEfQ7RRJVnWjWLz0qWnrOBZa7A7ucp620AOo3i1vnx4vcGQOUVrqP5EJLkkj3J
pmbNOpmHzC9P9Vy8wTo4Gx3uCwJNBGnimqUVKOZid+yAclZdcTXFMjfQseUcu4F7t6sRCvTHStx9
ppgOf6fLAm/QhmtCKj0igTTixKJpsO4jK7CTj/5AWItfBmAPoDhcSu46UJtzJBsv4PWEtWNgwbYM
XA22m4LOVxTbSPXwwUW9XSYbS56wHrk+VsuHMcd8dzKJoM+FhABCBvonClADLEqSCxl0pPcj/xv1
dXKellYz/OpSZkKnvSzGkdSOfVfX/ef9WKqnI5/rUwvsjgmRm/QLVERQLERgAOKypNpFFcOkJcLk
EQYL7MeDNrvadznLgSj2cgTYiKwQNGJgCsIu+v0T8UQO2zl3eRbjSr1yc29mmn5/VKRNfFnPH2Qt
HNRiWchmavpZJVwQQygWSpMRXY9odDVkvYYOcGZ+/vl407+aA2IXyaRpnkknG5CPG3LYZEWPYqdo
Y9H64fjX9b0JSVTaHj2S4AvWlL9Fgj2zMSeczJ8AhXbxlFI6HcPsdNuhmS0tp1DER9vMGBJViXcE
+G0IQfNIqtYy3lI13qLTw56Djs7/gS0bWSr5oKCjVxYpQzr8S6/QBt5MZX8/njhpCQ57dyC19lXf
hdBRGpaQ0ndpl48KGZ+vnUqYwgG6Q6yKoKSa30iBd+fjGMBdWMooslsf2zzXIpWfMet5E3HGkdxW
8L5NYhMR7HGtUWjjfE8xsQkGjViBcpfgiIBfNhG1ohpT3KPdrkIcSW/vxPUH0RU0T3wI7NEokGX1
WujMDvxTGA4gQXQW4iryV5WXC0n3tEqFfEAVXsQHcWeg9cF8eHyfn1LFHD/CCjr45+q+Zt5FKO+P
SfGzyAw0SZ8/dCIHIlO+FPm/dknqt7Y3CsEyKxPuM3XQl9JAwlInt4u18gKsn+ZC7kIoQZH8tnJv
SH39IFMmbgJv+HXDuZnIyUnwpcixLXuWVRAHkJl8e8qANHhXxa5Q3AnUwD9nVcJkqRhUrjYDZGZd
5iDspfpM4b1E83E2hVOEJenjV3TpFkObSxvt4dGECpaSY1PMk/w+eBUq+IC/I/FMzdMZnGJSvJlm
C7na1i8vLZCovTBMN28ChdLmF7NdZsU/iwMjLyZroURtb247aGUc86kl6WDPayk0Mriw7ix9rGzA
6sdeJor9ujmsdH2U6vu+TRsKI6Xrm3wt8YzrvAAuO2bMb1cHXO1CRG8UUSGBBAvLUNn3xsnf/n9R
bO+a2GHIZEV+LWeTveyONWw6RxVGCQTcADNukm/zIzsQt2spxxF76C7BOBT7rA2PGcnihL7GkkEk
kjjr6Pchl9ys0vbcYuselbjDDbohMIpQ0M6uH8SFOrh/ADRAXe7qRMq2scrgC+MlDxofIpfyY1Lj
jmQcXh9hGLP4nhjW2ZhKfNNjHNbmIKbZtB1lbkw9cz3xHmQEkqqHHY3ddqV5XJun6fVmhl912YnD
PeQG9XWYw3SrN62yU2es6eOkz9XJkBe4oUK5o+pJ/GH56WvTnRvHWQT3IvhD2CyXJLq2Ra0vJQ1q
SQ53Nt66mVLR3qi0LrLR+W/qGzL6yotmCfuKdYfF8sXTD6NxThZzvdQUWHSukdYES288D2EOcIsB
tvsCjsyEebG8/wfyhvY0IZiWqiNuHmV8khfr2cVVBNUODRsRypx6mDYlDnRUWfU/wh5eV+WwI1wQ
fKquiFxnGGnxblG0mVGq46fscxR5Ie4oKefJ/wJ1o5wwsBGzo7A3rOO7wlc2+aOvSU4EpPTTEsE3
1W5ZpQZBdUvErGGGz2K/DDeyP4P76MDPWg3TYClEQfdWdpSZ+MLHvIqfcqrsZpw6MPn10NnOQ5x2
a6s9jA9NdwjN0qJpYayvYd1UlAOc3R9nBsLt90Tg7ikeABHzSWgq4LbqDojefxcKcs2WFzAAxh74
7UF7JuB+oWKNoqOVsiwIUpfWejyLDw0IA31FtUMRi33rwdO/3GrZi+1G8mp0VUTD3vmy1bnC1gTf
fSgeb+114jYAA27vT7lnCri0ctrSj4ueyW7tN4EET3PaiMx/eRBL2xizFImeY00UH8Ku+zMtjrrQ
nFrQVu9OrVcW8DPSbWvlrysWhvajKKYQJNvbTTrEWDuyB/9hBsr3oN1debmOMIH4nYpWfnhH5F24
ZASfGxzPoiQJWg6YgoOsO15vRoDazk9LgUgbuTFEDvTuH72v3c4AG4IzA/MoVTwfBYEQCGtQ9nXM
5OAJ9l5Gwe/uXI4p8zS/iAdrsKUpyxzdRXPgJbfoeGNilS7a5oD8ZXJ+iqDZgxL1Y0hiO6qemXGH
C9Cxy12JifiaX8iaKj5UjgBFzNQX7TwoRw+6DPcNYVhBj0H5B9LmxCMkTQq+moGjpTd8x4B2yaZJ
CCiMMGrfx3ouwIk7qzFTCd/asEZj9tpsKnElNrPoXK7w1Z0nbTforrZUvW79IrInlVedv2t2o++/
/YTYGgtLbNnAlI7XIVtcTqAVbrOND4gcgMywKIRJrhwYzJstxtCfJ8F+umBBRccDfrUK9wz23RrN
xxVhR9HW3hY9OOWUWRGqPJlgETexn3U17bJy4BXyMy4Ifu7wAMjwymb+GPm8IMTtPtOZZnct+0FS
jMHOy4ezQq1FtzvBVMP74A19YsyH19vzY5AQRnqTRdVIF7nZYeORAJDZmXLLjmpvb9s5ANEMK8+5
TK0bLbwEjsNyxd7YNoMjbP3vURrPOhmPjX/kSnFdheYHfZ2SXFJhBakJKjX/l+iIAzaC8Qp0ChyB
Pa6MEWFEfCBzWI/kRvjHMZdr9INYkseiifIy7C+IttR+x/bvsdEFwuK3/PbwwkgXKibuGbku3/gE
X1lF0Iu+mc2il1DkLOei8/nIeh37lZtIPwXNyCS32Ya+iZfoQb7/y2yD4U0XVcx7mcoIjVrurRCj
LVHmhilW6/L80E8lc8xTCCuCF9cpiXenCOTyYvUKNyXta35ydV3q7TH10bndK0afIRy+vtOlnb4A
rPMgPaDU2XBULhdbpVfLFLYijJ1+NahvMNO4YGewE6hRQtNEnOTyKljTpAFHjWiQE4DhBJwJGljw
301++M6kWtORBG5tZTmgt698GydEYWH8e+79ZItjLeRpHLWFveGgFzl7EvEii6V4RdAYjHATkiz0
gAF7GTYsEIx8omOYEDfvZ7q/JY0MWqvPTggA8cmNm7gjhuLzQlavUKw++NuEYqvYm+v/2FWGWtvD
vWI3XtpcSd9nGtFgEEChszD4g/1H3SmMgfVQqgXtfD0enakRlQdC2OGakx2llw10TdHB226vhmm+
GOmCfgeqIKboQCo/76AuxvxOA4lNXi/zeHiLAlmtgky8W8AD5h3OgPqdwqQrnDK65K6vEKMq6z5J
F7C05cedeR4kxSmP/I9XtcKg3hHwlMJIXEC7H9Q5PJt9M9JBmSxHEhT+BnJV2Lbhc5t9JbyWryw1
ObEA92GrYS4XcCBXDbkIGlG/jCNGMgIzAHzSvGtrWP+mWoC3NLRhYt9LLYhkS2npSzAEQmm7nz7R
4Xc0Yu6H3yIOeku/92eHg8FzzwZqMTZ4FLibu4MMrTENz/joKGJyBaK8TdjksaQ5R+H1PFqSq4uI
NFyDlmN8lFt5dbQCWrNGToI6anOrV15N7bbxbYmxgcJQuYpjaLi1l3Fu7i3CaPAK/LOb+DilAlTr
NeBftLjPbwwXu9p9fUJuRw1Nb+5STC23L/LXn+NoEpZHc4H9mm5E+HkKH6Q6LfZ11ji5lm0Ma6D6
DbKTgDDQKJ2cytUy0Nwt6wfqFB4ss/6YSuJnGcUFeKCw1Ert1Xy/YXeUJBAXqbIZzGzrdOplMmUe
rwpGUqROraSHRWfNp0FqZZPcsBFFY4/fwzAye2ttOvURAlwF7jEhICarkbNRPVuu/f9/sDlRJWv/
xL+lSE/WCeG77tMLt4dXjg41cfVxi94sXh1JlSmF244Pyxi07VOAQmyBr7yd5OQjV7DrQ9iz1/i3
MArC7eIgNTrO9yJpVKdtN9AFoxfoJV9LOq33I9mcZKm/daOWPZc23jasxM1ezDpKoX8gST5396sj
3ExamoqkwNITlYh7j08Ro+QUmhgzR1sZEfk1PLYDZ6sV+MMKeBFq0DKK9alXwabaVzapnnaQtMzA
TSlSCH2N1J9RsRP2OPgcPnHg4b5EQWbi2osGCGMRHdRGYqQbvIlThFK7G7pREVfHy2tG9NlWAdh0
AuqCT+LKYM99UFju97TvSVHDupogYyiuZjFZnpFJRSeDEOW9z1s5Da1QieZBNrbSqxPoqeloLMDW
rknWQAG88fBX6IIjZ0Mq4/46ZEHfiTX2ymGRVyb1zRBvkym83n7uo3JnCFQUumldgWK5X9U9er+v
uhSsB6dAMOq1cdxy3HavqelVAgPYUd9HRmVInvnt4HErN/8bbjhVaWiLzeIMTHfo/TcGUp/QITmR
tc/JmnIjz6OkNiWlv4dq7A3beiUIjGtDdebF2vZKHKHY6yrV7yHfjQN5V/bICsq1nIBZkAmvzIEu
+ihmPyqZzOWK4bbGGxZd7FFF9tjpRNDo8Bphl6hFNnpj1YPlX8MeFMwfnuUZ29NzF62gqhQgkFA7
JixmDBOvZY3bNRMIYq0eNYWzH79tmhxY2MR6EaRH8SCOqpCVk55zUuZq02NYUBagDeoS6p/LZntP
SF4czl7eUcCmeZz7GqbjrDuffZjrmPnuC9SYEuf2Q2MW82XRqaAfICfoZC4lobMsbRgnXPYjkUFC
wsyOTRhCB/6/bVfltL2bSIkozRrGEybjA40z64CDzhMnBWvqWsluFwtDoXn9XD/Fi2hllUlhs9bH
CIx1ZTk8CIjgMFG12xKNRjpQaT7latA9CE3svVwaXR3e81hhWI6AAShWgZQrOhVqlUW6t3ihUO+a
I0qvLzQrhpG9N59x5ScQQbVCCnSOn1KCZrvqxdTCVuQPR4ZIi9CS2zTaFOhWIk8XdMzdfRa3lWLq
Su0NrU8BQ6ArSNMd8xu1ns1mbjLfen4o8Ri5SX5oMfBOQT2pXNpnQYb6V9z+jPJyW2W8+pNjuqNd
60qmCLM9+pLa/fKsIPK7pHMI0e/zVSTmkj2eme4U75VK6aeDWp/8ArGoT5WYrF1Ro/4Luo4S6hLs
LfK8KrZMOXoii80qXKGTT9I2xUuCNg/DKQKBjZrInYCxMXBwuEnpE7JCtn4JO568dX9tl0eFXT61
97zfxv/bayRI4qdqSVEWJCddv2m/20HeJ4UNNWMbSTYSnDX0SLwFI7oBlWBwV1BkFtfLHyyrlvXZ
6oPylZ1DmGe3NwNM6KfJKD/3KsOx7pQxWJ8xvfMDidhEgkm7uavsc0mqe8b6yLfr0Q2b4apMlC9U
nLm67b6gvBwU/Tluy1ry/H5UH5MbYGbI9ZAOcrE+E1VGo1p4l5K60auXEf0WcbVGtDVIxbVxOx5Z
CVn0AcaXgl0E3Fy4B1TUlBVt8TQQmoSueYn3lYJ93gSxs2nCEfhZArW6cg8TM/E2Tzy67uuirle+
xFXAnbaNX9MvYo+ZACZxFWw+tL1OxBwe78gDCW2+zJWzlFKq/P5QGUiwKydfVepd7fbUQMLOIc2B
KOKdRxcOfI4dZf11PERgXgAS8r0MFh4gANcHpO3PWMZx0u0H8ukXZ80g2oH0xtXmIGYwJXO0xJpE
VbgB+XJzbeYrQu4Abjd7nGqhhFOy9oLsgqQ7a29OP4O21XSSOsSCRioWkXCUvslBx3UigiIs0ygc
rpIy6WA+txJzS8el6OJXxJ8fwK0OTdf9Hi+ATBFWhmpTDv9EJ9QiS3a4yuqzQe7U0F9sszUbpn0J
kvQqeBhXcKD1D1734iOL7AiNlmMwJ1CUerQcSqVsTizfEiPkrv1Ve+o1dZw29IXOMHeTOHJwkO8h
i9QpcCYxkUQZwmxntwz8nd9cnzIjhxm4wksPCFdJBwIMSVgpOK6ri3t0U7oH+ZUfAH8dkyEvmlQR
oIqjQbAAbk8KBgFvlgnLeBF9FX0grAf05LIKH7a4vUti6zC47LJELVsFYNVRegIgm5Opk5GFgihE
CYu4zgyYfjvITkh5LdEq3RtgUnDnpHbTPy8MC7/sVkN3kfSi3iuvBX9VYaTmvtbdh9/4PxmJjmPK
vLrhLVc7c0dFBu80kEbTv4OXe+PNJezKFm4nVDuNwPr+ckrgX/ooGzO2dU61415XZvoFz3ME+FHm
OFSpaATqd/VvVFp63iEkuRpB91eTezkY3ot2ip3sEgmukGajkkI3bJFzLH+Fic841QsecApZ2T21
KaCzImXaiMg6l9/PVZbojsvePh+B4rFgBaW45BE7xFRDF9MKOcztCy+yGtRJ20jDWMmgiF+0KCTL
GXuzl0V1PE/v6J9Ndm3zdjCnjF+pYI/YNbwzAYfNMs3ZxQQ9aRIVoEE6FQzTo1qy7DvOhC1SzwdV
hu2k4VkuiTCjPVn21AYNqP0+JGaVsttY0hlCP50oCZBEcc6BhvkrVfMP7dTpco0B77wYV7b9f9sv
UND14KKp+lD4xujFw8EWurpdTHKjYBUx4jyNhQXQokHXb50KTcr6v4auNOdESkw8BylUaxKUSjC6
gr2Uv0yojMoqr3CPtN1Bi3gjXNksvFBajFOZdJNXL07grfPScCKrCqB5iMPseURKZig9R9BGMJkn
hCck8rn6PfhRXZrBtADWfkDd/dpcHramgvaD71/gilMBMgjz2vUaRltqybAmSxzfipcs8rWh2Y3S
VnmcQHReTaUedgNpmz2TR1mQVyLlVNEhqHyOR/uyFAzs1IZaURU7TnRidlH7iDE8YJdfgD6jZ9Fz
NJq8DpTqYhPH93SB1fbgWkwdOMDMSyTXGd4OzgEIFSBG5a+ZYxlTq8rn5XRbuil93+qlFJE2A4kZ
f7MXMog7U7h0u3QtFfusoVrN2EMCFoqO2GsP/Jdch8/aobBCCa1HyeDSyKwHnPWga1vxgjjh/iqE
Mz/GLYE2Owl2iTu0IToG29Z/QHyPy6zVeLn/vRYeZE37GrhP/Yb3nBxYQOmg1eC34DNGf5nPPxy6
Zv6ZEOX4CYP9LIxVqDKAC/tQJTRNvmTE+DjrEx79n5GEZTQorMDZqCHbKQGKR0xrEOkiVNpfgsvU
dHp6kK7QSTLA36LVCtefy2Hx4Bt8+Dmxrhtb+vlv3AvqDOuNtD+a0ejHjEziZWiBsUqLqhirGPoj
cVp1g5Bcay8poHQuzDKXJJsX3O9pAfCcdUaf651dSJ0GUihwGFQWC/90F0s3ZjxNNXBsKSR3Lpbq
g7UddjOY7fS4lRvBKSjUtod6K0YE+cE3XtUB25bHAqxAKfDAkon900sjTJzamVqYTVJir/9rhIcv
f9C6HVMP/pzq4weSl5CUAGfNzN0dVONqiYvI/oT/gdFJ77XTdJPu9LL+tQlp0tJub6pBsBen6J+b
KuvXqTBMtr384t5TZzeWwkSxTrtH5Zm/0Oa0TBnkuVrDrzsqHpOxXhEzaJtO6rZf55EjbDKwHl7A
I+JP27P9hsYPmR7TI6MxqjpfYqEM6f3uhjZuzcGwC0CViTG/xGEvF9rYO/gF5eZJHi0FCNjTdP4W
xgpco0viw4HtB6vhgniWlJgsM7DrdNQTrxzv4ALu6RUklaohuiE/9Fb5drhFt3WcWMEO23UOhv4O
TM8AFa+o4+IoRV3kYl3NlpNkDg7HgTJOl5QJaGAGLInOt+eVSuc2gafjEAcWiUAoQU2vsBD6SuIZ
k2bOpZHfrHtXud9E5ZNu/PgOJbhxJO4XKvsoZPog1nE2qZnOakjd6z8m2LelHwitDvq59iadhSpC
PTs+o2lOhAoYTnWcVuvbTHmB9OyKUBvbEAi39f806AZ6tfeufdxEfhglAchXaQR+N1ASJIMmSCWj
/Mq2kFLbo6mbLV0pYsrLqsyLmJXh0pRIVHBIs+8uJLeHrEMxcpPG/abkgMR+/noHZGtCcXKJlAa2
or7Rjem+KLFp3OlW2NZi/Dj7hvVndfJPz5AXh6NNGLegrOXDuDaOBAPIzJX2sOA2PE9BR4A5KkNF
E0mN4SA0z9oWPKl/O3BdS60MXF+RaPeRAS0HB1ts5f9tAEaTeyenrOIDsCQWXwsrI2JFUnMCBDD+
MratmdQnQI62TJcCvgz3t5vQFNpg8ugsmYaAZ0O4FegbvvRRLRbBewvsMIuMIwR+ThGr+0D5Ty9H
x5N0JRPUOR6l5Lpsyf7NmR/eI954PffvjZxHgS215HJIwzY5Gb76CDg2djN3UhoVFouzWIjc7ILC
ZYQYTCqPqnIxFaK4umHLZVCW4/FGYH1sQuD1of+rKGvZmJPeeNVmH/k3nrdhDzueQYwdnF5sqoXT
w9hShZuaTvS8wv1HtXzlLY2/exk6ZPysYLBy6Z0YlzYkBqlXEUWfmpdjVsd0wG7sQDCHwAyHQ5G7
42ysJUOVl1kcHsQXYEK+htEalbeFD6w6PokUQnpyDQ4QsbZ/QhqAgmZagH+DXbRQ2S7ZD2sDi+64
KQ8L+x13z1LNQVub54GtLLLUhTlOolVkw8qf67M2tmVSizj5m6CtfL7PbT9ziQg5INCxBh+LaxZO
jUEDtQ+1up5xYHkAeNAiWC2pfhCzvqdXaCYeKr7HXfg27W+BK05H/GG1l1XOo30VjPRmcLaSxjfu
dzPrn2vvzncNbMX6Eku/RDCGFCz/zFXvQFG0iTdutLIIMz5J76UApP7hmH2uKzGtQ2QE1Qx7EQrL
sdMDPOeb25/WBOTaUX6N4z1FgDs8iwOEmkwisafiuyaLWeHP90wVRT5jfIv0/s03oRItmFj6UWS9
izpBLPTlqw7ad9cp4AaQp5/21Xu7lUHyuEdsIZgW/oP9fh59QWRW+9D+o/WHaWrXErCiF9QVW5ke
rDCNjWTj6PJGlzDoZw0F3wtiHiypMv0gqnIZ2yD63GyPZNoEsCYCJhIwhdPv979nlopcsXYMs4VF
2Bdo8f+bFHgbMWrNKVMQ8phK4EmxByeWS61L7unm6A4ZRPUtKCOJePG0gMw0dtUXAl9Z6zpkQPuh
66k/auTX3S0SsOXmEVfRIqnUdCn48+rxTEAt9WsZKvilAHtK5HL9CaK05HLMKQPjSMYos4Gpn8rv
5Y1BNvqAfCjlRgAMAXBeeekSI8HYNB9/LXEjvTAT2hHdKupPf5LBoHeXecKgUEAYqhx/TqcPVQwg
gi/ho/cJpbmZP1cD8H6gzPny9WtZ8r9i3DCmp+fkkJTVllV87mrhkWccUH7pDQD/96NRgkI04bxi
bblV5M2A0YY60BhS0p4qVlFCNdyuZAo1d53Vyg7fxru1yQ+3YO89LH4JYkwioAWK/hocScsL/wGD
F+HmdK9HEhbZuhwdsZfbm+P4mpK6WaIxT7zDnBf9EdDxXCKJi5B9S8dep8lsohcD7xgPFvrK2ltL
Y3PM54h0Y0Knx2JnTLLZItHqFo9JoTo208lDT7/KF0tRREnMJ1wa5iwF6TSUujJvyV5DzpclsD08
ljocMACOI2OVT7UiIGSUw6bMz1o1fUbPIOSqou9CFBWhnehp3guLipA3OB5donQQChh9AGW8B0qN
BIcLTbNM3RIUPUlHWxp5/x/da/tYEAarkQ/02uIfYlmlIcgUuqQ/F+QKM0C2SuxdqhUd00lDFt1/
KRXn8eQd5ySs6tR+S0cOXXLoli7mO4hTAIRAjRpPodXozVHO3xZYMMa/BEGxaSh7AG0LA6gqi7EO
k81EjNCt2X6rKsDnypLoYe/Ytm0amtgpfvzfL0kGH6/b/ZfR8B+dC1lyxZoqIY/A8WbS2MEdREjb
cRDFhGxzxcAahUg5Xm1PSg7iS4+ZUxCFpL371G4gaGUdDAPIj34lYdOM6/IxKFi27i8Zo6cPLAyy
sjeUdS+qXk+YI67Tecc5uEYQdpC4+fXKOmd++ICI/JJBoYV94Q5bJzSmJmvjrCoiKGuwXqu2eyNF
SZwoU3H5WiOOtfQR4Yvagal4cuRDZ6D3ilWdd9Wh1qoritUXhUXnHV+GWAq1X0d4QIO5gAJ522DA
nwDX+D/NHAB7LSqKz3G48JDoOLWVPCRaN6ftet3Adir6L08ySlE5H0TqS8T7wAUAug+JpOz9l+CK
isZN8a2GQBS1HCImVO+StEsnAWNsd96JWe8zmziziQdHyrB6w8wiocE93/rOCJHU8vt/4UfHfgm7
IkPUwJQEAsSY3bnRfcSvw/0J21/k1RDQifaxpBgWRPsYMiUmJkq8e+xfDTbqFS6rVxmyX9pZi976
OrBcD8zThUuAuiR9T/Hq0h6pYVuBd819hnfQsZvMqF2YFIkgyj/z8AtmxfYpnAHRzKHy9W3hIlfL
FvyCYBgVdq4eC7AH/vWpV3WSHjJBRGDhPrVYT9iS+sHbrnmgLPFObSvjFrm3kAWaAgNdThRKZpfZ
/ykXd/8noV5ALPDYEhhtw8p39XCxpVcaQ9QgLGdQ5nUoKEDPFvzMxmzdFPSBEOG+hIi90e0uQgHx
rivWbega1G7omM3QT5XwfJDwegMbbZ7ZcoM5ycvS/9+po17CTFPTJkDuyNCaRY6iOcEmMmm35b6a
InCMfxoFKfbiFn920znBKLNUq61gaUJGRjfBXJCa7a33PUlUw1NuD4QjnpkngMSKEKxZJ7XHQFvR
hiTKj1NItH6H/1OI2YN6OknqEnamI9v6p2019oNj5W6CATMgQ1BpuneSuLcurMC1I7zYlvZbsP0T
DzKL0aQ/XfcABAnvlxXWwHaKhaR4CGjGckh5c7aZZe7Dobmav4DINZtfJLEotHdgMuaIaUhuRr+q
9LPtcHJdw3y0ri/HBVOllN/Tx1lPJCE5H5NNXiUqMt+H7290/S9S/4eX6RVUJ0+12hnlQf7PoH+e
hYUorSzFWyHzvIp5nig5gZLPFBQcmufqT0BayVqHiVVdRkl03v7HcssALNzDutFtIkALVD3OnN9A
h5S3OBZ2v/lAKYsc0XFvWOe8ht/mDwEgAdIhXt/g4qa5LpCURX8mDfYmrni/RJF97BQA7paxY7BR
qKRAkb9elxLLX+z8BbaMp4oCWTxgawujKd6EbzBYGEspp9Jaj1eWK8UBb4F9SPO6g77rf5UQuQnF
m7acjLO7n5UhBHqcfnBgY85ayCR5wUHp8i7k7giNBzmUyRk55Nnso6wPFi8EayivCrfJaozu7ly2
wSPBIxwaMNrDX3AmnfV2MCvHPJxXl2wKI3x2yWQRZ+oxT2Dgnk4A+zPrRAZz47PktqmG6jIxPT+0
8nDlVYZbuq8ufPBpeuuhzI6GWOWm2t3QpO+AgtXorc1X/XsFbdRMhHPNggzD3ZKCjp6gjdUq+Dno
gReA8srDsVoxb0oujYEnOZi3XFCApQ865RH1C5Qsl3ONX3CRHeP5NeIyPhiqM5/bke4t1mtU7Fse
ARfFsRYEiwzgQRVh6cKSiu0HrJvv7VrtPnIoPPEv0lK6WSM/t013Ytht+Ob2VPKowYopaJitojRv
M1kPg5yKFLq94KbDDd6ZStTrIppeER2nHSF7To5Tsbh7vTSHDmOr2E+XaRs4Xxzjo8/8hdII49ks
Xb+zApdINy9eNC76+JwgcBg96XL9aBwkMAzHm0U9PPwD4OFIoOKjRfzUfSmrkBYrXie+iw2BOQQC
9RLzB4NWDMfQ4hpLj4A+CwoSC56Pve4/wV3GWLoUDjGbtVBYAQkflaFkp9zR2C0dHQm8tSWqJV+G
tw8+s1MjRU7urQO8C7dnCmYLe5AzNQ1c2GfUnVeOInl/pelfDFyyyJb3bmwYPewQLYmCgeHfoC/s
xeQLF4ZWf5WV7oHABlbnqRYLbnzRmhx2jM5wM4VkdAG/8AOvAEsy9OVjKbg1AMXuCW4o09KekIFX
eDjyQvHv8JAf3B6/cc6ILY6EMUorJiwDgVxOcgXnhZsYUKZGV6hdm25dDjZOhFuPbFCI6bFZsQoK
dYe8/6iMfTTvgkAVUIvW734Ea7rgp4+uwnIBcpsvFdKDjsL1okWS4Als8URVJs48wVPqsu/xVZvt
wBkt13b6v2UtvpJyfQ4K6yr+GEd+31VeMtc/icrd6NdmiP6igk3/+T4y+x0mflkh0bHWaBwxCAtB
a4EWkm09hYmdIch83ZKPaWZ0CgZ34ATeSxoz/9idIWpfWcLYuGa1RsKscyILrYhxA7ckZfJJdaKg
qNMi/zN8hZukibWhBO/pjEsPHVWrIqUbVf6m1xJ4xEfElGhFmAdFL2SXYLjIOgzzmEo3Mulmzbxo
Qv8zQeVFMhUCGTbUUlEKvdjKcINY/bg1B1bUg0ByWVB3TjKRzT4pQSI+Xz0YY2A61lZ3HZEv/ej5
GZwk9OgWjAyKYWku48fE1Q9T1VnWO0JbuvSwT/zPBXIyWwxwg6Ywu0P+qFQrV5WMEO77gwMcamHz
aAW8vIyHOemF4B/wbV0VSlFZqKYNA9KjpqT1uWn1BLytZRQM3a0sZxCIUhc7Dd7yISZk2V8X027m
xGctRNcDfR0FFSbvViRFyInDlgDsSDzMDJevz9u90R7FjEWfTtQFlQpGdS8Tknh6sRBfWNs3ttyI
oDzAZWCdmWYj3hfWyM4eIv4gXiWNFpyGMsGe96CK4fx855hhHkAjp+B0Uoe9L3QpDxwB/O2tB8tZ
yXgLvur6Lt0pDphTz/NCRM34I7kZ6AFinmhoBftLvCA/mxsgbIF8cWxpoVUfqF+DugV73Jd3tqKH
luMcXAGcRJGgX9yiIK0MG7RRsa44NH9VQONNr3f/+Lj1+4EtoEgUpNQpm5i4UQIjgqq1R8q+kYpS
YoEh9pW93HtT/QPXOsfY2Js7NcmOXXvF65MK24LfT70esMkcIQj7zZYB2NPPqGZzgXJoRPoVB/XG
VVdu2kJlOo/Q25zkMVUTklQclHUt6O5sOtHZ/KtbyWftM2SuHaKf30EHabB36nP26DpDc5BSDhr5
uC0Q1VO2DsukpnD+IQKInXM8tCbG9B2d8+To5hTfLL2hBANUK32hFt4ka/DXwE2Yj6pkIiPdr3c4
bfWvEo+u6wtAu2xO4COjfT8jn7jRXcYTb8e+i90ONfzV7F3k/L5WNG1t0DnGcYAur4jQSFL9lirn
Tb86EXNNBPYkrkzoNWQ/zHENjmiy/z+1di8Dq69EYA9xRsNpg0E9+SpkTaFvMk09LOpCAwFbwtrO
W1/+tey6aV1PHDI5Mfb2T0hiZr1ym7cxZymra4BZJH60V0LzwsyGhz4x77SSdEY2plOk76geafNw
EmtonowbjWTl1glesc4/4R+VGMosJhobJIAtbfR4vrwjucbNuWhDt2MUilMdq0FuC3OD/P3e3YSx
Q7eZpZuiUrQTOM0yIwh/CxHWsbvlx0Eje/+nEEMuS2ZAnSNBZfe/EKEDGzszEKtkzkxIWeLxYgHl
I+pL/NJPLQ8SmcapYNR1BVU8FOhz45bkwuBj7uga9XvX0zJwW5m0jxCpvHwW+vxoV48C4m9dQ3vt
Lwdpffm19FAfR/9maoZ/tejNemrBlsJ5TokM4hI8rco7V+BHi2dnoJzp8qY7LK91pdnurLr75LDo
JZ66rCEBiL3271RcWng7GFH/5akF9P9xUTzjZYZPz6QUtRRqCcZu+vp/lWCqZl6ugikdbDEU+K1g
PGAYDA8YM3Z+5CHvpYA5s7RrcCUSuWmu40lCXU6bLF+uhd+phmYEjG62DrKymMTMBXS0i+PUQ5Px
/kerfBMPr2O/6awfGeINewem4kZMBfVH/RPY0YpLLAn38N+C/DyC+2LsHdTeBByJrY524CGeKI3c
HnsBuqUFFUehkEMAxrOgzKZTZyTiU5jQ2mzzw9jiHup/f5rjfndXWGR7F3KqLCMQBIK06uTShWwn
kLYccSd5gpq3oCRpfgWVzBLB0YQMXIK8VcfV5HC/haPcbla/SF2YLrMpy1HZbZdZ1i9rbYUFlJQA
FOBcMWYE3E4B7RaVX934sknsNHRJPRvyZB7aaKUz5uqFDiuVUmQ5mf7lrTE28uO/QP4XXuP2Fjoa
CyVc/euqFhr4WNApui8gwTWZLbmX0yyl0aXxjwpr3LUgzfdOkgk4HzyxQh/MZx1VXoDheq/x1TEp
4kmRgqZhZmAMCjHor6myqsvn6MoxPba8gm6d+iXBO534pl3fGV+A7HDejLPvj17yMM/3j4r+54FT
iuKFFjFPT9BHYNcwTxdi8e59VymVTiMAS/ku0rrDHpIjZfgwev4HLwmcH6x7TJKzx204wq/CWe6e
PYPSixqUSgg0Uo3j4Kc+orePTpbh8t8WoDfUVn8XPCXp75t8aeRDtl4IaFWTC4fSVdbO3f6vLVsq
b2sxq4ATHr6/era6JfrDBvkzqi+vMO1oImJOkRDHF17wUFRKcbZVBghJ+ai1xJ0u8L1OwdHHUGH0
Rp+x8138nGkmU2QmbwF3pxF+97HICgZM3lpw2/YfryqPjWr/mexNdOK3x+4mJM5IqMK8K5jUBWZE
MyHFfI2NuD2pwKvquE0EpKN8JHOEFT91G6kAyv71Xz/Uo+jCzvLYRuV1qAIQIioEiLdCxtCIwoBe
ChBtjC479SHLkuU947J6HHCGX1VzScyv7b1HxaRkGTO0Z3qKXN6RSb7g/kSRyYBowoxtNuCiXcWj
cqH3RcoKyllVDOeuMTWmj/Eebj0s266ARZlcp2YkUwt16vFe2Oq5nXTtoPgNPsQ25dDXrI3CT0fz
wPDJQ8Q8QV/3d5LTSvdeHydoXaF2uVjcnTfEk7XY1Qt+RzZUfqN3OAp1VikVLmOqFaJ4+fG/ADdc
X0ghgTX29k546MGjpzo0Fgb7WUIlejKiH6N1PBehUWUdOBseZllUFSnfylDDjNuTBaeXOSFPjkWJ
bT9ooP8xeJR+RZIfqsXM0pNREeb0ZSzEsoK4inxKOPgU/hQ7l+oUf9YA5yXtG0wcQFpUgqfe7GRd
ZfapMRl6I1lqIi03bKVZz0BJoQgJgPSBJ5Rxp/OR7CJ26x38I+y5QggqWLTqDKKKsSrgPdVxRcMg
L/Gm0QisqV0fO/Crub99SmuApxYGiYGkUQ31Zjy36Ysr+XXbr0fgTqUuHmNRGNkQSTBNrYCj6Yq3
IZCGvNz8DKDghSZAe4vFt3EwSW1AAp5xr2TpCV+V2/z+5Y5RbI0gQhM4MZ1B3AtGDs+J3z2UegeB
RzZNJXHj7Vsx7gCmc0uPFBdn+rDePkhLknh4DkZD4PW3YmH0vyn4ebjgkzZnBAYBo9VdWLexQpsp
gU7h8mq++2miL9n+FMfgLoJToaS7BFOrdVp2PNd0kD2rltKfli1YJoeyFcZf64goG8fylMq/S252
bXj+fo1POPaqr8XXL61EJ/UVnf3uBKzRcZnwihi+ZVF3dn2SwOA+5DZhR8OMav3Myj81PP6faxRH
oho5gjEC+FGLl99Jg/n9YUxFhzVjGUixvRmuK6FpesIE3Mqi/OFxPH6jb8mKvdgumUxRMZ2dhlmd
/9Aeh0lhQOaAq09sr/8HV3wtCuwDt0lnl3MmZitansTaVi68HVedIdalmhDB8w6cLEQx0mHJKiO7
DRR0j88VR4rvPJPNsi1tF7Qi9xVSTmJSu0VnP5Gpk7wqIbnYx51cUQpmXQVbCoJauS2FpLOa9KKY
DIdrgrYIZU+lstqdLSKzbiAatSigeQeJHa0L521kc1kP1NL/5MDtuE8h56GwCON6m4dgWfIHcBAf
xjosjonTdfRl5FjljUW1ZkN00a7BEenjI9CCE8Z7QM6yJ6diJo2XefekasGGnXuS13GWlv5Uv7z0
BhrZggZIJ9w8qiOms61lfdfZufU5efBxWxYcwcmgFoaR7aNQjwaKbhIeWdCMlZRmgCvO/UY9dqWE
7sin9MDHXWPM9RMiWk+3XkvFpG0Tt70keTZzRlyfAaDvJ+PZzGbpANaZXiycOqIAxUTWKYHgh+8B
sqHnxfuRWEuRB0WCNAe/1yenZTJTk5coRiB0mdj/g5GTxRlEgl+rjrvFx2560Taftj/JfXLO1mbX
06v1L+VAUnhdGPDAorYiZU9cTCYUk3lxIV86qjhVuL35WB6vVhYl9BNULbVbqdYh9dIEBqcPH80G
K46YkXHPFcBCQA10S/I4EbGdhJ2W4UAElKKX7Lyh+sAjRCprgcI6dUZYOIEeTWc4/LYHZLfpgyHO
vn7F1AZLjDpppjjqzrkSjZOi+o0Exf6IyhWyzTwD56mWrYUZqmk1sEySecr9GEwzuNjudOYiNxM6
mmZP7XGDdtn96jL++5u3D3NQzR1TNx4yIXEgiyENaoNtRwwpB74ifdzXB/DeP6EUcxeZikSKVMDS
9GpB2AfFl8V8X85v8oiR1oRCXnCMgHPnUBKich97A56IYhIFXmFY7E717W5z/Q/T7Z8nw6ZasqvW
45GjIVRfmvf2A0Gz1p3Rnb6wZ+P74orjQgV6Iuvu5Ap9DiXme47fGzw6cejlfsGGSBj2vNMgGfm1
aLhLobtOXlRFscsSQDqHeoZk8SFBd9pLlMcCxSUxmWU2K+LUw0C4ChtldZXs8YW7uU0PvFZBB1dx
Exbl0HWyo89YPWOaxXgMMJ44KmQq+RTiMjbuOOidx1WG4O8ndX0E24o/sNQUPj1izlb5YF3KDXke
q9VIHPAtirbBAQEJABaQX2hOL9r39CRUEx8gmB46CprzDLRfzVoIYbD81mkOngaalC+rwYUnPFzv
qNeYXs8N+2iM99pRyAA0VACl6UJ6VKURnjC3ZHdT7rw/kOCpO1k+nCbx49ltRWDgt02Pgz3ScC4L
n+KMLWg8H0fTRXIrp5iOCcegk98TvAnewJmuzFZNPkJimHCyuAzCrjeFVLEvFpfql9hDNFbFu9EX
MJNatAvZho+qccEaskduTg82n1jPRng5DYrNukaiT3axI65iFkq63F3KFZ9ttCu/NmRAPfP6SW9x
wvE6NeTASg+0AlZUpvn/rjzMyXchzT3Ge/maxS/vllAyaZymQ/AorXLGjRw5HcoISRmvOM99/3nF
S/qx/9vttriGL1HK7X/bKYn7Zmq8nD3CwpJi89+5DF/vUIfos4sPpzXeA7kuzFRgZ1j4164+3W6S
nRluQjNkyn/1fegeFE02vvS8lGYYoB1C19MRZmKQTe3hLb3a4SRrY6TdYcxUySbhsCJDu7TBn2cr
1qmIJfcGXUOel/C2XIX8EF8zvyifs99Ds6trcZBj+e1qDZCOOEGcttpTfdgtBncrywXDylpVuiyZ
4uMQ2DYB+p3w643U9/RiiwF4fUC4fDn8S3p7/LWZDugdqYxsYLnlBsmnGpVZ3xg1isoSi6po5xWa
T+tQQtDgpuGOw1shMqaX5QfdnutIbvyu8dNAAJqSlsZnajj9WsHQtEOixY+NPRo/8+BB8o4iiYZw
zSkIFN+eUDNCWy7chwBcmvjAb+KftplYdSbjBAaGWja4RDd5hNorL/e9bTpkrl3ZycLputhu5pBU
shyTLRRnKxZ+JAPE9yufE/D7R7c1uQcxj5P4d48iJzufHecoqSbfOHVmwZEbLaT3iBs1nKKfbk1w
IUSoedS5Pz2IX5N2754g6dZsieMxhDNYu7ASIDDigtcthOoUP2BprI6kMN20j3VU//ltmCTI0Jqt
eEHVQ7LY1kb/JlV8BruwnTDWdmvWprXcCKFUD22QBMWwvblAWc6Junaww6wHr0WSFobZ8/IHX8G3
BTVh7iD44S1NByqMMR0nEPdhOCQLiP1P6mpfTSCWDGPZ3MqKGevW03Sfsgyx68LHrVpuL2wjW3DE
4jh4QuKe73bfvSpBQDEbW/yiUH1IBNvPyGub0i4WowZGQ3WTKpTN7/4Poy9j37m/6yuaf4NqenID
fIK47+uKnOcABcVjOuvcrh/Wu3DyRvPmLeQPOfgXB9E4BnbV9IkEFBlYqkUZe9WGXi2oJ40zRgLo
q+RYbzDIauToTfuZ4WSYhb5m4WVwyloh4R74IwucVmsyW2YvNxvpET6qPUHinU9FgxO0V9khBcGl
LCiGwVuNsnTqCasxhoo6gP+JyJXbbyXtQr5/QsKkC2l36F17XEA/hLroAfvSvjWawZgtC7sCTeHP
GfonWhv1KUmwZZkg+GrtNjkjGEvbHRqLRvnDXE7I+gTS3LKAL6wKNvC5e0UhHVS0lLPq9Me8xASE
vi5n9wqM9Ir3JJvQ+/oewp0nJJZHBiG7PIFK5mRxyfUy2zDdCNeNOGDkA3jeMsHwhPcrhGgWMvjQ
oYCzQhDCwSYjB1FL2WCozXYHo/l6UVV5Ck8gQO/H8LwBkP4Y6Nb2YY5+CEn+XCqOdBwbfy23+lUl
22nHG35t0V3+IpJYrAu6b9P8LCd3IQH1oQ8MB9BFxCn45hz1qiWjFL6rp+ifI1tQh2FwTqyODOIq
15w9O/4PnShx1E3r3/FWdYwAr2yxc4kFzXka4/wXyIHL83+DbbX3RmUT0pBf3b7YPrB5nmwHCILw
WG59IBiIR2La1NuTiiwTGh8ouV7DeKcgjUxz7NKOTYp+tbDkAhmhAeZ0t9jEYGClSf+Z3lVPf5xg
esBSLprrKWWuRx44VKrosCEeFJs/UawmC86red4jAqptRxTMjOZ8SEiMNh25SIxZ0r1DuiSOhFDD
j9eegUzbOaKWwz4I2ujoOq2bnWTNKIBVgpM7IODirzY4K49B6LGyYAPGOTmFXGW9VOZ8+3/kZKqX
OgwqZ1CDQWDJk/saSWoyd/fuh8weHeXvjyNsYg4bTnniuIAKY6cc13nfwkkMNXjf80EdUpC92WYj
47DqK23AfiCZeH0kL7JACKBCtTqn1jqt1dgGFgqNSaAQG5HnuXjt7y7ZwdfGTzQ0ZORhtVNivXng
Ez69aglY9w2h4qk/3vrAW7cwPXHBJVG48ArNwNDCBvH7IVD5ZeyMCmYgBnxFdPJWNpX5LE2U7AJv
695KeZh+bKHKUzofFikoijN0e4OxyXY924z/uLBV50s9rxGvV9Dgyok+lQcx+u0PT6gwtow1dVmj
GvUMyQkCE1epR6L2hRJVO/+MXm0D1r9uHCcq/2KX9murdVRvhazc3UnDxMswgTruawvrAcxqNIa0
Eby6wPRjaj01aujrvoa1UtRYQ/aWky2AIjMfDpVRG105uKYvJnLyt56HFZHm827c61QNip4bE1mo
sPDOcv8nNsM1CdNcXMVgA/Wt39wePHzXuoPl3S52Wbm4RvPSaOKufkNEclq/pu+tBDZJKx4QGUcd
z35HkOvYhGAF/yjWIxyx6C2NFvZx5yyA68iE9QCpWumGGf0xs6vYwjQj21B1i9X35c/7paBVZGzP
XLvqaTg2aWrU/ZHC4X/8eNZ98iHWLgYLNS+qVo4rLZDc9K+REaAFo1rklE8+x+03/Jtdzsx00Pti
Dd192ugs5mFnA7POvtRcn4P5aYKWYfQh99oPRxMm2cVF+BpQVbiY0/NEN4iSsI5UN6XUavmlXgL6
+VhGXgN/ZUoJ93O+tl3hgxgqjEksYFThN7rg35drIlxBoXmhprM3tOc6N62bMPzpGSIRHfpe9JSY
NlihYC/meezo+1RMdd76ke9jM0PMFH4ZDYYML8g5My6DiKDqsFMFer0AZvI48ucBOZxisTi9Bmpt
uwUuMoOWvVyeWQ5eZChlw+p175p71FLZQJOLKV2v8nb1rWIcyqRaekjTtD3sKs9X8GdpBsorf/dJ
N6pXf3F0qxgMIFpxaGCS33kzGGSvpTk7824UOjzlF3+2cYjYFlNzWv6nJusixZcIOyi1Lvd1Fb5v
gKof8SHA2hsHUsXm9xWoNYjbL2U3xsPZQROwNYqByf9aYHRR3tED7nywg2tzwMNfxeJePMNx+gQ4
B5XBAc+8cew8Zkv1Rdute/1ja1QtdW/AFU4DfY/v7syiIU+FgJPO0k98vGabkE24mYtcwFvi0Mtm
EIL6ggWpOTY43lcq7nLoRiOJgZH1wv0v7Z2OFXUCNVHYyUT0E7ZVkOA/D6lmDckG8mhXcRLrzCJl
8YJxkjY3U0fkZaLQUNbqAoVz6RTwFvNqYxuo7YKakQEZc755N/lnfmlIK70f+aQHFfxLLANgnhU1
nZ9tv6YRaBFd5C70j1GDeCLwXRjitWRSd5lz8JuX7yjMChRyp74lioCFJV4sVInoY6FzNDHbmad7
g50Qm6pJH5rgddmyyKCTLWeOI9a9OcYQ/kW0y1EhP6WoW9lVsCyI+Zl69ftZwWygIxL3qKjNqTFf
9dHu0rDsNpYr3gyEHFA3KPKA6ZwzULfxLgZHxOMDBq3aMoThYimQ+TM14l6Y66GjGPjBcpu38BUb
8ky+Ukp1o3x7ytv+EZ5K5pP0C+n/q23DmLDGPS6PWtPF4t2YdqIuaEqZZKyNRozYeeKZXDdlcsk8
Y23OBejKTZGv45YqmCgN0PALnoRlAGZEmxNT9ElS0DfAet8c3CWhtdIlV83VmtjYy9lQUlSshA26
uvanHbiwDNQ2N3psLXPh5TLtTwgSItCq8H/nq7DS9qnn2b6kz2+jH7BhNZRaFQVlkQK6femUy/9w
vYkNXTNRPTIjFzH98qblZjJiexdY42F3upuaChmnJjYx+WNPqDy4FZacNziSZWifE+jFQId2Ac5v
HZf4rjTmxNeE1FGRBm0MQPjpERjeZ6Baks14Vu3G7a/YrftKQT/02bWA7brk1Owcm66g9GLFynTN
VtcSXQrdeS6fnK/QrbPBDo2fC1XDsFAI0q7RZ235FQ8dZn3+CXMfqrxr/Xpr4/yysCTshuyLMgKf
XW8B13goTCwwQjfckHYKe5B6h/rO6Rh4wM17A2KcjvqJt3V04uHOJ0nrXz9wpKDgsStdIB2qhOlz
PQ37eY1Nag+3YZjEp67OHEAzsdoGgt/6yWrGG112YE4FF83zn3tni4c5Qs2x4NVfq0/Ii75NZcdT
3lYi/sS6ZLgiC1LeZcM9V1joBkVEPgozFXnNcwDudQrncMzrlZv4FPvVc9mK3VgQlS1fqkVyfssG
yHzUk90gMYt4NgAtz4d3fxyWa6/1xvYMxy+GhWEinHA4TT7FA3dOjy1U0q/1ZxNOGouaEGC/ta6h
73FyjwqU7ZFiGMwtbUXLwuW5LGgC+1G6LIrDhvXIevjzmWcrbo4woBqSZaal+Ts5o1+5MuKJFF6w
P/5eIeZ5cSsGFmcUZ5H9buhtagcjU7BPoSC1Bn1FZbH/er/ryD65nDUDLqTf5h37ZGSYFrTtHXR8
hrz4YOCXskg8K5TgHntDhbt86euE4XJKz65QbIl9YzI9PaZLPUDzwC5Nx+bxQO94S5QyGiPd9UHw
TuqI+QI0WmC+2C6IliJHc5jobi+vTSV+6arzfVkwT4w61HzAcFYSfEqQE2Udy5puIhcQ05FzFwwd
v77GKQLVfSe2ujSJVfTw8bRC7xlgqOZArqHZovICrJQwkleFRNCDdlfRu+q6B2w/BIk5v3YViFZw
d5lWJj4u1nJi0p7z46Ic5jhUQa0zj7UvhM+z7VUE3Gp3olWBSFX/3eL3zFEWp2P/uKua4xLwsaZr
dtSjW5/bB7KOe1iMlvq+LkohvoESlbsYTyLvnW8nDrR4nI7Ax3MV0IZ8Wsl66fPAeiy/u3HFt1uS
8FbO9VoUZbgmKW36M0CAGV5L04dbJEgfePKX2GHgGTAIQqJwsCVZ9jf7yUaoIq/VG3hskUUv97f9
lnosFzFMMoPa0793DVsgd55BZpk5aHLWNAMkObHFwRlEumb3Rp4NSEGz7bH50PW/osotIce6D6mP
I0BquqN2ZgquyTQuom+l805VTClrJgTLeje4da+stL5O4C1zsaw4zwmWgIkl1nhrCygn77bSHJgU
agKUyvclTfwknOBh41eap0OwC+cdAiTUbe4gGjfZhomIcw+fMfOP6igr3YXKgfOnAS71ecbY3+xg
RpmN2e6Kyv212gNObFq7OPXns2pgIDf3rCdKoiyQJukkzbO3OQkipdqb++RuHtfVXqic9RARSyD+
vYU8HV8NXL5P/Nz+Vxvzie6ofCHacoN3sjrAogZQgpdBspGJqdwLPGTD0tk3lb0i/m+lIUWQUIMN
lHImVBswoe9HTBN6gKahE6Hhf555/lHVSTiUSQSotoPdhJcRGX+vouS726okp0+4I9sbdZhR/Z/D
N2EtlBDq16sJGXPzM/LNhJa7P2VebUbHcfQJ0KS+uUaL7RQpBtGuInOf+5CRJc3tgxBtx9r7kf8x
F9d2civQ7v4zKouiAIam342JgHBgEX89Zn+UqKyCgofeQ9IlH0giu0MABe6AXhzYq6Uzu1s8k3xk
e6kIBqJmzy07hb9NnaQKP3P755V9PL2EKL4MweLfwjWYsghyA5Hx3QkBKzdGTZroISLNGc4Ih0dl
YmxhO5Aeg7MTyrcKWBctbW8yet4X6ThJBAv6Lf/nqLgQPpY70SGoLw+YfWKZj2h8UiEjf64qWgvs
s+QaUnuFzpA7dRy4bsnnss2hetFVYU7weaN0/0uXechOD1tXAvDRm1fN3iSnKljOc4xv8zDF+UKm
cuuhT3gqAksgtpod166uTw9AqLwHelIXb9SrbFBCD4AX1KEenxcTPtESvgdgXPds+IDbGNIvg8Xe
9Epr6yCxRwwpVlzVnjZZA4qKjoEiEj7FoWxwDfrlyOUw3x9zf6tp09Wvap6S+X24kHCo4UhZgWJz
HdVVGWi/2TVQVttKJtw4qKKgk3rA/Meqllk6LC+UIYY5ywFyB2C9nL8u2b08+RH3HW4BZGHxFi3M
Se90ydoYshhMjkECLqjYke822VpjLB8HHQqN/pWoeuSTI8QjBF1WRl7o0YdnIJBGS70XkwJtWdHw
PKDebZg5FS5EXOdG3N6luJbWRLrWMrtFdLI+bOX7lO0edwRhIdwTUjrblXF6T9ypE2UwKv4E4m/4
02mevAh5vzlTAJHBygQGGq8PP49EbUgpneRQ1do4ofNeklGvoUPHn5p2SwQCWLUJ7qzuqqNH1UVw
hSPsnafWzeJ1ln6vdd+nuOlmQ73j5LbLWGCyO7NKANNOw+oiX5QhuS82m//phPyAPGBzn1dCuTBm
5qRMSYFU+YYsq31GtEACjYoKVuhTimezg/5AiEZnaonVOF3A2BQ6bdFC+bmvXT2irVTmxG3AHH3S
Qh0dXKfVocgSWruipZ0St9xBj1tNfC6f0IwtgWZUju3tCuOY/qu8iv39oqDFCWDJUGFdWtB84f2I
q9qVZ0o9FbnY/o8S8XRVkr3EkH1jmU+z/+Gh4NNn5QobbrcFnz6sZfKn8CzLhJNtsolglPBYFBDe
lDWIyPiKY+eCcSjtBcdamFpcXshdg9IO7Hq7Zefh62D3sfz37yum51PF28D+MUzdo9ZimiNizt3p
Ltnl5KEShKlPdT1qu8AyA6ig/L3FGOadzIuRSYKG8icn5BPpOzuOIGMc1AYdmCdYLTkg/QxJeWcl
HkYtIkhpRm7TZp2AiLgwn+jMifRtyMsLf7/jpH+fayHjfAY/Zeu1u8AjyQU6YgBINt44UuffqCCl
+2f+m8nXoUP3oEB/qJvUm/nSyjQyrRy51AtF0Dt28HI//kA9jFqLaNJYW4wMnpFo9M2e1/XVr29J
tzX08Zl/45xKU4YoM+SozIb9WOIcW3UKf7hkWj6kqGczrMb9d4NOfXSJIanPjCNzwFIP5dnraN+I
Yns2y9kOXUxiBM7T510O8zK50yV2Y6+Ap++o7/GLaiMnJKrzDTx9UISeb1kAl6cJEqM0x36+8r2d
pjZNvOXT4T55FobnyvS/JDPeQFVvNJ+zqVq33Rbnd2opuiGa1GbwV52ZbN0T1CSlT5ASP55VOrju
vRO4BlXdMPOBvtnkz+wttZW2X3ALTSOWMF6jTkn7mFR+LY+3Un4jfD4FCH4cUl99Ticfn3nxQ7oh
LrBT/YfD7KklLKEB5a2W1oxtDM8xGxR1RlcHXo04VOm+C7LxE+UEiFT4bseLyrXzblEDhwLgL2PB
0SXSGpimzGxREJRjjovUs/4kZzpUYKRijpGvA0BUzgjEkpFMNzo0gDxab89DcnAGe32XQo4w4FQi
OFKHqxtB9by+Zd1n/pbnSmTEj0Whad6qhInL2nU86DyPs73l5RDoOj6zCFocDzXT3jlOgvW768Wa
uOimEWPNp34cQjpIBtdgea4BhrMbbI7DZWy+G30ZgNQ0v2K/eFijGsBcCA2XkpMqLWLlmK6Sihd9
NDD5TLAFSQelXcO9EbdjhHeMKgYCdcZoBfG7cPEAxvG+4zq+FGwHqs98/BGddhDct7bCoqrNxLUc
U08Nw/wc79cB0IM1WTwFIFhkfRBmesgZjqzH5Cidl0YImVADtQVBNmLUE+trM6p4Bb2GruShVYZ6
HEdP1up366u/CQde+c1hiDC+iz9cogXpmHprjFsIZCqHMLU/iqQ3frG85PkjvRPsEbN7GEyCHZbu
Ju8IQplE/7knDm80RnNKtoGc8u1AYgwpNUjpS0HNJ+lg2i3BaSDop3lMfeyXVMhUzJsX2d3H8gHk
lpuNhc7XnRarUAgYk5VTGRUJCyLZM0NJup8CaHYO+OLNwbYAL2w4XctRHAJV2BLINuMrfchidoZ1
yPOTXC1C7g4DIP7tvrYVob6BxcpKxD2gIv3nPWrA7stFmRadcTPZdnvnks5sdZkxtEKVo/0FbFFI
UgptqvU3leXQifYeGZ35QkIACkDlNAEeVJVxoLw4Kf6g9r8/aVAY73NlORPj3vG5dUezjgbWlQc4
T93THIgj+2FQmNCmM3t4DTO6egjdSw2H2nUGynlLElMh9Z64MTqMye/RnYBCOwAbEp+Z7tfB20pf
0owJ5GsEs52ZtJwHZGQ9KDPpdoVSJRYY3rmjveBHWIyxb4872rKqsIXeIvffz74kSWG/ALdddaTL
ytW5Y9tun0O4s2r1PssOu+80VXlA1vZj0y4ilyVat/MG0kmBAgtTrwsQmuFK+wT+fiJSaV5v/uRC
W9p3bMAnKtUxMNhvM4QaYtrd6XigYlwvANt9H8e92f/MIcMCSKwNf0K6cH+yG9iZQKmJ963Ty+On
r03bXOcEha7GI7aNQCJc60XwRyaTUvzlzU4VUyH0s5Y9F9mD1wEm697jIZdUx3hnbgZ3EHYJEl8z
k1wvXE9a0dA2NTMCMIJklamBQtYKcLU+ove+LuMmPBdBhDCEbrsi7Ud2DHwL1KqzsobVeCptyvrS
zrm+FTSwPaokrjHlyVKSph24JRk26MmPE2w7OG0fMNQz/c9VIFlyD598UETAfG0MXJ6Z0nL12+5p
HOdDVs2Q2STmk/CdzoZv5mPHE7crKqYNNgvWU3WPLMOoa1ZzLB74gj/aMarnS4rL+Tcj44SOcxof
yOg/VQvEUWUQY19ctKKle25EsarzuXEtkZuoY3/n9uzRmuDmvV31E5FRPcqwUDi8o33ecqwl06mu
OFvLFI3PRyFarg+we7jgh+4tlItTVgMR+2l6X6M5yBn8VZJmktycX75tbFEjv5dgFsvst5S+ojWg
RIeUuNzsCEyi8zcfrxwXcJ2+TINfSnFA80yg3K6V8qJ0efAzS36gjRkxMzNvC1Hy67Owi7KceYds
IOYxdyckr6OQu0LztvP0VKjVklP9jybpV07qzVB+p6IpPkg3dS2XPoQM20DkcyUpq3FR3lvnwZcT
A7M17hBg7FB/xX5df17dZQKCPqiWJXams8Y0mZu1xtSjYViJBecprFF+c/xLkRILbpYUyF7QgYoI
yC7dUySHFwDyXw659OQvx+/NdD/EZbCT/TfE2KxD0JtfztOCt0UzN2oKxa/o7BzcdhPSboW5j+w9
sq/zQf8ZFozY0qiK7LNCw8Y9PCFCjPAoryZV7ZKu9s5LCqeHP+XQJCsjFSbeY6vQpAI4iUKcffxT
kTeUvy9OxfT5TOLxE7zZ8BiCeyaekmkoAGEPQF+mc1aofH2n7uSA/0yUYJJt7aPteNN4HpkICN2l
8rCRxPqazCa3VivlqJ3Lw9cirVHx4KAW9DtPbI+YzHplliVeOlwI/1eSVEWoy48hQBR1HKaTT1lK
1DVkjO+3n541I1+ifLcCC5pgyyNdv7wUerM3dv6QbtDpGg8o1+UvCQ5yPfcnd73gQvh++Ch3Re7H
dMUlHIpjqsSDIdtPNvfhvhZD2RnSD9uBu37N2TWaJ9ZKpZEWRUdiHYfB9qaWd6P9yXF9e03EjUGm
vdmbpTZdpTrtVZjnhoIvBqE0VAyvYkiG3yL1GcJ7aD4+R7s9PwJXQOtR6NsxmRgnT7zuIrggIL1N
JdCV40d2zcLRfskpFVkmUr8/p3ZyJxqzAxQhAU2xOMnWEulz/NuxX8Ske7pua/QoAbwxsoO2vFSn
Zcs7nF4fYWwg9fIUejzpHGbScmZMuroQD1gDzAaSHXtQ4LZrt/OQt0WztbdICntK+clpb1wY0PHH
qx3on2KPWiQ5QZkHDRPkMu4z7S+b00lAxS30y5YRtw8GVVeIqQZDhJAo6ArA84va3dNTkC1ubCn1
M/yed6jDSiG13Lj38E7qu+s/Q7LYORLqEbbB7ZwqokFp20+UcV/e33kEyXDVco30o8vhvD9E0nxE
aNf/hn/GfKUhn+pwZaBz8LU7pTFdwtPCy6d2P4rVFPkZGClzMYHYxwO4QjgbL1oEuPJfjQ94wmVV
4PvyM5TP73BrdSsEzJS9Ere/ZjHvcJ6YxOJ35x3AkW4W8yrKnsp9fuwd2+e0QUeYWXVqjIQVtC8K
28t1jVlgnuLqDfuQl/YEE0WafQolh9E8TXxQm0WqTqJBUyPdlZP9LCd36gYnKXejeJRgbtCc7yOr
mc5rsAcDOBko5MTKmguK2PmVjGwHL8M7A9kkBXaAV+8IdjnSsN/WZj1faQOAtVbFyLd3nm573Gpw
vN5hYLM9LlQQP3dcnvO9iZPohZjic+279o5n9nHaDWE2fvjC0q76hK8x+wDf5Vvpbl7wHbr9fWXn
uS1JE4LAC2SPQpkHy++t/ZCpo4anBQGO5S9smKequdRxoVt+W4uV/Znt6h+ic6V2pmDyQAuNQ4+M
8p+kL5r+2tx+6Csr/UB8ZQ/9WuUjdl8NFBhGPcP/xPBffFnnI3Yx6i5gw5CnlYv1na05frcDIu8c
xt25BD8EKO9czxbVBQsHEo8QRljPkRJ/hRnTTQKzXQ65KVPZ/MCqhaObYUP/i/OMWbiWJToLYWQP
avDxHoLaPqgtY9MSnaS4lUBZ9p18/KuMmDfDu3/2sjkXHOEs4fSJZBiFamY+r8YGkPVfsMjdAaZ0
S4MLEohwRbO2v7NiQFEi904tt6MdaYye9XWB3Q2cfrj9HCOKo4IY/YALY2xMcyA+Dz+5NpIXiBPO
WWHwr7pcpNcuUORjrVucV/5BYrN/62tNss9CYKKHiVACeY2BZTvxRsZQPg9ix57betwQM1xEZ2BL
9kVoY7hv2tzrmCTTYgaVw7J12koGxhYoZy/TiWK4cQ+RDwMpSRipM4vTUoNPqaXc76hq+DI3L8rE
tqzQNp3N/oNEYTxcxRoqHElk9b0/1/bzuvosMZ5jYZQ3dikCXtXi3AhggUSUVrKtfyvYizuPs5cp
SyqHh3SO/WwznmU5E9npRc0wqUNApDTS5z/phYdaupJ3ncNYHuiUylypABRyog8TC+X1CExj/3CH
FGKccMZYg/W8bTOu+KBxSVZ1ff233n8x2ryTy/++0EuAqY7+v7vJTsDBrxq0/P5xYF0dl2lOyo9T
JHgsGSc7ilkDRFjuzldDzk9Wz/Kp5ha94AMnITSxC0xQyFEqH/AZTnrStallYO0xGKP7/YcUUdIa
zzZc7B3YyOFE1P2kzmub1Djuk27gHOWa9mK78Y7LFGovd10gNwQwbC/JNj8F/MTm/oakvY4MBvUq
hhVlrqjwww34uRLzw+0LmqZJsc3tk2b+FUiDF04tVJS0iKHh9F4OjVP5djExMO6mIltMVVSJEXHz
qcLZBf9lCYEHfLf3Y3WNTcpApb5fcZlHiKmD2weNol7p9cs26TG+t1xwLceY3pi0rbQoUVv+ngVy
NmjKXMIB8Sh9cw0+MCOcmWOj62zFv6XDkMCLIeDPpiaZ1ttp4xs35tH1u9TX6xUimVqkCjfcdC7o
I5QKSQdmRbE9TfI2txECKkNa7ur6G0Nq4t3WTgCYw9s6/zFFmAOlj96OTX/jQPOLZZvay+VRe1f8
tLBGXyCK1mCUasFWId+KP2/a3IwrJDkUuuGSfm9yrxtlFdWnOCa5hjsAhgozrDTWzCJgQc8FAnnL
3Oim+D42PMvv2viEK74ZxKq2OkYmEZkNUOrVstMi8X0bp4lusD2X08fxXGGQK4N3zAP7X+JiQGEE
XO+1UfBIW+bbdOJN1uYEFot66Kxe+Zz0+VGbcCSQpcg+D+tv3zomZx9wPRU1qJD1KJIKJFD9ogFk
nt8dSAl7bKsSFd2a83RBrQsteKQfpBEAR9FX8mSXmXtruJ93t9UJ042m1KcT8meKko1Xz7jjFKZ+
vWZ4v2SylRceRxD2IqILRpevFj+fVNrj2kwzJC8ksHBxkPh8iFetoDrgg+EIgBZwAHp+AHICAEy8
WK5FGO8PznZfxgzuwHWj7M8BhnL9704Q9hwZMExA2c6UdTPrRgwHUSo4uQsMn2j8TKHkq50ERzCz
wdCpf/Ofy9vx2ao9ypugXnG6Nfg9K54V18V1Xtes/e1heTerV1t7L2GYYsqWbpoavjPrKaxRiD6E
tVK89yZA5sjd3Pd2C5O64XxEiaeixKfwET/CqEhvyfnmID9qmP9eEmlOXaJl8+cFT1RV844V4nmm
WoWqjsccJ5rb/CY1jRuiBBgY6RPLXiMX4Uhs10X7C4a+oagV+FieKPVwu2KlHBOm4YQ857VtuIIW
Gy2DiHo/UYw6HVsVnD1u/uXBd0HUrMgYG7i3Pd4psQ2Iu7bF38TIB1vYNrhmGx3ADb7aOmUKBVL6
MYwTBMHFTsVtrDAiQCjXfKjyLb4Ig7cZpkYig4R52+UDfqi9b7HcIN3ZYoOu0UZVsuikFAuKZMk8
SamHiv/HT8fre3my/lnooORLZiR+h3O3o5h3eAD80USsA2lvOS51FJHSaZ8Ny6YNMMRbvX4xOO/y
BhyRvJxGvBcXhKjbRbVFGmLMhOxZ4QIZRIFhGl9QaN6Nmh2N3yxM6tGPf57i+9gaLTDgzzIczPlQ
W6e8GwhuIAvC3n7GEMZWtqCQoB3oe9qc+y5+tUF2ch4VCspkyTeIOw4Mc9CMBBb3nQ/PI0iNntIx
ALq73gRQVjtUtRElLk61YYtm8tkzBPlNzDBloxi05kzx08WtrGCpHuw0/GoOMrNSextxkp3RKW+/
eDWT6hc9xP/VmdZYVU4bX7NM9kwKeJn/lbDSNpdeiOes2LydGxCRGWwidOyxbwsFETzhK3bSQ/9W
hcnnehENUOhj71kbBkaoebCtM5rPnW/8wrqt+oANy+VAnqciCxzAf94MiiakXNvqpathV2y2I1xQ
AbzoF8lPCdgzIQiN27U8mR1nvdWOcJdXjt8pAo8EQgRBk+YhWK8cW8UsHFjo9QIbuspdS7LEXEBG
JWx9KtxFjeFNlhZISXi4tjryqMtKkB2UeIduGLNr4fwxyMBYZrRzd2y5Pl0Cfb8OaxKk1BF7eIED
ZIJMzs9l33AanJsLDnGAUsm1ridULYkjjATppNjh0zF4EuKq1fcoBdeb5x2FL5/xkK2iAyoaic8F
RToMT5o2sB42zw1+az4Ie7j3GfR6AnAGbwCQB6CJGvqXJ3zt7mMsRGNy/TC8V80B1dV53U99cLXq
uEFJqxghgVHnS++o3fAon0yKGlgw656r8tm0wXg+cg0UAPxR8FbzxBvfYe+KrQCafRLlTHQJIru6
xmmqo/pRK9BCPW3bM2d239DkAjjcIc12nX0PCGBcMxRBesxHNj4xKdijY9iPS0VvDKNIflt4YqU3
nB18HYG5LNc/nN6PqTy5kLEcZkrytvu8A6Dri7D4d+RHv1r+KWn0vT4GqejFUVcpJ6AMRCTbswTn
zCojbgJTDLlsv4kJbkYm96Zkx8m238ICmWOx8aO/Nh48EWrSLSRQQytZoq58qilgjEUB1EN9RTBF
46Es3zBdQMVaHLS7fikAJaRhXWyDUCcn/czNXzGMy35N2BNxkxNJAjxtPhuS/JBPlL+bGKqaX4ak
B6sgEnUwk+DoBNn9+smBCxl6AcEK2xU9oHBNMSE0h1j5/0HgZpRu9J2DtJ3jcbKQnuotFDIzSjQQ
EsXIRTlsFNoAoTC1fQv+40feLHsNVok9TYa2HRoZFNFix+3TM7PcD2SAmJih2z0E/ypqaMfRXq9o
Y8vf3Cez5vB6vCEUQltVEExHeC16Q0nkhw8cV7HhO57/Jbca5Nrsu3O9n2aOmltWLGyr0dd99Onl
eIlrQ6AUDFYFOU+FbiOuV5WLJeIwqVdhWKJNOm/FExKgwipCVcmLdvhJ5rzJWLjJVcwLdvHunF9E
GWyZbCYvcts+1U1xYf9nJDc0E1yi8MPDAkiVFVaci9wrrKK1nbaplRfZFmI9wPo4DMiFDgIXKvrC
A0vynHbYtrJVACMz7mLUZXoHjCVV60JPegYUm8wB6SqCglBXlVQZ7KQRRIYZCBjx6wCSCJmEgAif
L2m4OOheJH6VNYQy7Vu5ZRzAhgxGHrHQFpWV40B44xzKPf2GOvC1178KrCfBVw0ajhlAjbhttQ9e
m8R8pEJZyPweQSjJ28XkZMm/9VZGanYiTU+4yx5aEXfthd0epRjhNEwjnz+Fr8ouFUt9odG8LWjo
uDf9RA3lEl6YvGaAwn67XBdpTW4HUPIxcvzM3wJKmD4zs6FafhYUAE3J1bgoG/EROxyNKEJY9B8Y
p/B8DakqDh5169F3QOegnE7osAgzyx7aV5xc1idpZ5vySu8VtCGm5LNFUbnHT/fDgeZ3Orv3IZmE
DJCJkRosUqWmV0hLoU2B8+y4dSOkG4c4eqVLU3zyE55rttiR1TyiDw1nLBxEketdbcHf25uI2f7B
npbh3SPCq66ItadXkNHuLVy/rHAy7SEOIwO15OU/HnoDROFMeD0f1qvqMpDcqZEIaU2KnNvOZXVg
MBwLhIal7KF87XAaZyZt/EFHbv7ZVPXzz5CHREgtl4bZ+JT7083ZXWDxS21FBMBoNbmUMVD4aKBr
g9JM9uKOdbAtsmRmsu+Kclg5IITZ/cqm6rDG8C+zngGcoHUbN8zXpeBc7foH7fjJ5dwWdFPxmlVS
CutfKcJwkBRePSx3L0LvnDXOI/1q/Kie1Wq/SCMbOMTicND51pYnDMUQVqquXxd8sM4sFODgAWZr
UTBm4+bdfulO+IzlqwDCur2J0ntZRBAU2BHHLwiaR6sk9/IstbdyPH3mMcqQ4okO8IkYE9xh1uKH
6Q1hbgEj4rkZulRhom3bsm/num7Cl937li70YlBa827V3KxNtJnY9/WbktnKfmB54SQIUyMzrF2P
llehOHxutlSUHPkIGgPXtSVmJM62JyiJUn66YnyOk/YaQAAcircT4+FPHcTZfC4dGRsl4oBippcd
ebGTHT9dIQ8zeJnd1yYT+jN6db6C5vrfxIImd8oXWRpaklkfadopZynet1uMSI+qPOUp0gH4IFVA
XmxY1a7t5h4H63ys8Je01F07i39DXYfypabi/MBmBPit/wrWcGRobHT+EYnTuYWSm635kYmgnuTr
QuizfB/bz3498A9NjE/45b1bTF/g2OJuldYaZyqlUz4G9IrRHGy3bwx4KeZIOPfVPDbZOr65gqCz
f4UPIkmfjxZsNnqfOohl6NICQjXhNoqORWhxfDneRzebEPbT54bj1fknh2kxbcbKZ6Tu5sZ5hQ/z
tT3mJDnhiuaPsfFXtu5+8DuV3O0M5UQBYZ+elLYQap2w6fu0IFCPft6qwazkffRJugrTucVX7sFs
V4fXGRxCV0mShn16JX3McUz86L2gGAt1Ix6qcHYwL+wse+NO9mshV7RCWlLNRnzkFz9vjmF21NvU
/7hxbNODWwI3nWFcI46TDMSOi1YAMNjujJh3mImxP1+NcL8o8ViHsv4mrALfip1tW7jW2cqaUv1n
d3STRFvOmpGqXVVnN4xsYPxVbHU4+H/rKPTTwH7BQRMIRKUG3SwZxnhcx2VnZ8y6W9fPLN1IqnmI
SgWKn/72d7WqlltmVsIY9KsHckvJTG6gQesPvHcs1V/TTQJOIWpPeNn9NEmzJo7OVLDR1d43Nuj0
lrtR/8gdBcP77B0rh8yys2ZbIfyeDq8EBH9Ehf551Au5On0rNi7ErcJVPxB2xXqcqHJNFdDQjvKY
c7dK3fvycPE+7kvyroNZ/8koqEhwxcStY/Gw5xkueix099/sdkFrvDZ2mN2NQh4lBafDHNUX+yIB
U4kDq/4wVdCqmGgMPBfWtkUFesMc8cEIOoBWOuJa/Ou2I299aiT8q03bxnEUnMo4LUaxfY4J8mvN
qyRxbsN4gY+26E8POhpAl6PEaESe4jgf8RtTywuw65Bj0urcln1m05p1W2s98ki/+gBbT11rTRxa
lMP2+zmjDD4zSRtaF3oGyxaCi8VRwPIRaF5isJYV/3MpmMWcYVKCwmpRu+7UmUwM7ECKmg59a8Nx
HJST0NpHqFo4kN5jNa7MCBY783r/ee0RUfI7v5fe8pmpTXU2ycaJIVHFdg6cYi5aXcrgSZyv45fE
ZiWEG+q1Tg8Zf3ULAV9paQnRdahTMMt+8l8bcFtPhBtP3ZbsHtDNlBd68DyfbbNxCpVokJJLhqnd
lTsCtwKL+sT5c+pA2ZASP6Wb+dIlBT4g7Q5euRFF0VGBAUJP44lMil8wEynvHQg+EVEpS/HJqWUP
KSNgjUM38RlNAHjWKriRm1s5ZJaI9ep4L2nAxJbMIWoTy8/+REiUxlIOsGtLdeVSH0XdL8wZqKrY
SwETylkPP3/4eY6pWxupBW5zg61APfBb00hQ0J1UQcFRrSi1JVsrLIr3tyyIthqogS1tlrfFfl7Z
KEb59mIzTeGDj8oslOXwjPF/JISANQcqmcLc19kuNQpWsHqZvi4aMnjY0VU7QLIN5YA4r3RbXrGV
XfzoSn1ei3VLXqsasubG0HvxLc3hhlcX2VGtkj6kY/GZ+tMc4QG3O1Dg6dUYVCSKxIk0fJeIlC8a
7Cc4/2EByNzML34vAN5tCsUtlySbVo+nqW9v5Zf56siifhKAYW+kkCDDseqqkFxmINdO7nVhiMVh
+GFoZZxjnupormBBXvxzkZiHnRLpxJjMGG5b9rGLGSy4DBI6+aTbmM2D35Z8cpPMHYU2PHxsSVo8
dyhZKhiGYJfoq1X+RagmvTxMpv3R7Jlt5iAUc+oe2zKn4qmH3btYPWhWpHIsXlkKScE8Ss7TCDKe
KnqrvPH9SX7eomOmf184knvUwzFxPyxOWq6CoykzgHMCh/T982zv76I22i7nV1wRktPuqgzMU9fO
evuz5cIWWqo3z3HeAIevH/UynJQ6ROrk36ZisEz+ErlO1BK45riJiBoLl9MDD4c3t1MWwPOuDA27
KwmX2I3vzQ0BKYuTQELoCduatRdRdeCRHQ5/QAJdEOv+kMcbhExCYg3dO3YwIV3SKLNAaXhAzhGM
YCF9HL5YuIbvlAQUc2ECSiNfma3ixPQm3IcN0dmaQqM1HvviULDUGmYdtleAeeJBJNs8qpbZYWwF
7+JHiplayyySOAb7LvQYn3kXMe1ShBnx26ba7c3oo51WPIF7jWj3IHQQqWLSET0M8/aMIqM69+yW
26UeQtOCwzkoI1/D5qNROVRtnOz5EJ4Rd7R8sGL1Zin0MyHwJWzPGER4Gl7iF8xdCaWvmf598vo0
n833jSIYgU9BBP3EM7HJa45X5gfLNc3BdaOEqMqGYprjUoWXdUzusYNJzCE/f/mNPGogeeZteVvj
j4SB/F415aVhkx5aO1HeX3Zn4Ocrg60n9/hTqDT7AB9c/E3MdViiUm/hbNboF/6ax1IuM/SnFWOI
aa8khAgrFHyMKg1EQBxbKxb/Ds1iUtqDZQOn+24XZlwpuiLZuuQU9ZshBZfH98Cz/6eSCRDORUw7
upvhm95K2iuktBMTm4p8v87aWlKzp5ekWw9Oh//ploG2aAxBnHzjOHmTNDcwkud0nSiBZN1YOb/z
L5jskWvMEmzT/a8NgVPE5ZV1YyXwZjVPvTRfmpT5n42AemTTmQjD2O17172xuTUxsP/cjzWfxxi2
F/C6/bZlNqe3XCgjvjDYSREseT89zs5lm/TeDbWit/dVwhM1DwpIir0w0oYUCvbJYqiNH0GeHDIK
/CsB4EldroEYAcSdKfoK7k9SOTv1crLiRi8ysy4KsgOHl9zAPNatFteUTXV5a4zYstmbcf5UiHmz
D230oqt6o19VDUSp9dlSmvgIWjWm53G9el7GM9kD4WLpjYmauR3C/TwS9pytB1LnuynQNvSRjgpy
bHZt+iKi7vZMS3hq6LMfkYfYOGRKZHdQSDMrFNdq3PpwG1IqrfZhzrZ55utIzfnBW5ls+VfLbCyY
Z4w/bVXHVSs/uyK/NQH8GDD2sL9k7H5ki5PRzNKu3CC1rZmD2/lWQOz85vcVSdSJ5l4KcuBDolMa
0whXc7UH8ZX9RRQzNjlZVYxn02BaA+JSewXittY32gsSi+9E7fUQkgSddNX43BGVtgbQs9ld3ltB
FHC7UnZ+jOStqex63/qWC0UasIubXZSKrxlIBTi8kmrWcxUNP1lbUBeAorQet95hAToV3wT7R/Y7
VijWTqmSR7FYZdjGoMlziQsKi664x3KDpaBBfk5GuspVGkJS17L3x5nRJ1j2XBEIlY4jCM6iZ+yp
0iw6yKMi5IiNIcIl43N+EyBw0pBEteBCtfs6P+PiurFzgbQsxDsP/jKurLwEHM8mHt+oOtLmMeL/
hKDob+Ne+NHQQc1h+JoukBb0Yc2ZLI2utnNtUxUBEWv7eKXDb4zXrKr6ejzXLuOpYWpKxp3w3uUK
tyd1pwxGrnlv1Cfc7w2r53uhF/mwROl5FPaVbb1yw0wpq3Fc8KGUgcQMyPzIohy7n+N0o9Vnq1lS
wC+PSCW5TVI6h9FPrxKwy1tepE/fWA8M74AWvMptS54aeGcHuav5rpjGBDitPIhEjVDbtsOvqIbW
/7S/ed1KsLhSyqnKshZL1RIuvRxTPKPq/v7c840Wc7DwF4huz4VhT1oInfhPWXUNLtXxnIjg9qFQ
G2WG5N+P1CzRf9/7aiuOIyNfgSur+wSpVYMTNuHTb9DVwE24L4B9whJUTIlv/Q/3trbUVJClm1+2
1JncJbfuykephL0hJZGueiobeCEbud51ziHOg5BE5cF+rIbyvVovGYxjMVB4670bRKSOgeuvpr9b
fNCOft2ysVbkXTsGme1xCzmuIxuOp0KN2uTJdO5ohJPtBVbQ9g7ItBpWqA2vXmoD8JyPN+7Jlb9V
X8+jVrYKD+cXIOwZxlwWKRY8P04/kEwwnyGUJR8iRkItubeIPzM9E4qN8kwIhvaM6L+JEGXi17e/
CyzMNswo0i0bEULUCcitUPnyvK9dFxKjaswBvcRddOwNNuwp8w3VC6hTO58F7wv/STIRPjKJgxfB
RWO+Rs0RUgNr48pVGAUjwITr3lQvywUCUj4TQpX6+00czGKdj6iaGB9CeroBlfJ8rWVL0NglTdsC
CFapLkt26yE3LBEpAbvd+jILky7kaWcLVYC9wGMo/l9eLO9mphBDHB6kL4uBKaaHCjcIETYvUiVF
q7UlmeuExVQCeTjY+RjCVPpK61S5749jr0kmjsIkns5xoPQ7Z7BYu36U5EBdQVuZM7g1M2aiauBj
0KMMUPQO7vyRmC1NwEnSXNVIuyqJysQDvQ6QfA555JbryQKYjuVgiatXrXFtDgMJPpKRWrASf2+A
TjYc+iliLBaiQt631TYxbwI/463XdHlL2EAX2napsm/GAf8y9rqiTicM8+jAQG6tYD27+G0dhzbb
F4lzvNiB3ukcMapYkDabwDsAjXA8V5ju9Wy9gzg15WCHNWqmy3yE+VZh6zY2zoygQr70eqGc0nrY
Dw4dhrg6UhjcFIbbN8I0u1d3GALsncjNOsiC/LmHD6DDE1EjYL+zgjmeVDXeT/wimlsAEUC579PB
DlhxjUsLgCpLgVawGETyJ8H6DowSVwp95CLQVYjlnFkFeiOgTXaff7W3skg9L+TsVvPhGo0OFppL
RYrBrwkuPyca/7Vh8SdlPJ4sMiVbUvgL/fFS5BYrtRvo0cPyT0ICVaEiI2n8M46kKIDS7ujwANy5
BzubNkPxH3t3wXuEGqh4VHGlhetXId1PwA9LuxAlXmGPhIrzwVH39w6tmxuWCYiYsvSedX/YAAXT
aViwc+Wd/PwUL1r8UNzF+TY6ds8b4oCPt1s3wxti5kADM85ldD3TId+Cgo02XLwiyx281nldbUkt
uPx2WalLU8MZBA9+Cvh4EX+ECE0VfQ6XTiBXHaYnynLJpB5LIuw5y1Zd27VVjFNbAR62mc7T598F
iOjz5+QZ1/UV5H2ShRHUl7MdPlCU0avZDzzxSCUTDES3OovsLQsz0bMl/R0993SSOcv+FlPa9hMO
XzCPjC7MJroZ4Hk3v4MjrbxBCSc8CgLIDYhfvZ7wQgOr7zWSPj6nOxPLuEmqZ7B1jd+AMg1hh04k
EUkHkSFgbmcPFq7wbpdeAoyhig1lgWrkC7rGj3qaZS83SeS+ys6Km77Aro5h+QxHDgUkj9iCjl1H
vJdTMBMfN3d1xnBuHRCv5lBQZeoik+2g5lswaXifZyZIDiy8MzEtsWRS274Ulu1T476Slz/Cqoia
fYDYaWkutVfXEbnaJ4JDGPAntQGCxaIu+zn1w4ch/as1646fIymix1FGP/wnELVNLYANotNQCp6d
Wa0XKVXtDpxTEkrGuszaZdWbGoCLAJPeyyqb2h6nOc8oBrQDnYcrgqRmBdwh9EBhD432o990XdHz
jwyRIEHR1WT1WW8ZiEAo0GkSm/gSJHqe0RmbhsgZQHEjwb/vIe8vMvrW+NlkZGM8VG4dQpcNhcWw
/30tbIRjEzA2zTp2RdfZw6zfbew2jpjvNG0LrrcCGaUafrDVOTXLf+W1LZ+Ue1/vILg/+QlRcdcn
yXIrjMKV1KT2r4lYOrFVDjnUdVQcE0wo+h57wbhes+VOAWVHNClINS9Ld4CcGbOPJpPHYr5UH74Z
fyj1utroijahqYHiq9wrDQRfPkRqhhfQCU4bjJerzGX/zFMfnQTSTGYQ8JGqmngQr/dRi1pwjUrL
aaAhu8IxRmjEAYlYJTjc5VcsCi740uomT41Vh1l8DUhUFyhqou1s249q3EbenLwn3NgdRPLUMyxE
7SA51e+y1VHT927tyh3B6JHRj3Dhml0NrtO/pCedKkKVyC8GxwzHbuAvXL8S8MrAnY8jG1OnK50H
dj4JBbmmYbHiW5A4FYu25VEe8/Y3vT3vUARHKxOem2OyJCY2qdPF8xfxKSwPk6gwSZdEl7qmsB7Q
WOlcvMxjpFi3Pt8DC5rvrDqAeWYT+nriIhAZ9K5Zc5GziD2hYwV0W6ZiBj2MxWh/KmBoIjwGLlrx
G6tISz/RrQRyRYEewpvO3wFzVuxnAJxn2sDKS+U52D3MrCLibyCtXq5MJgNV/r0CPEpCC05xzE4P
qoIo/yLrY53uZiabJJ+R+xoymxFAiG8n/7vD35DY3M6h8X63kfeqXcfEGBqGMqtFbtkpl75GKO7a
WXx2kwlnURjxxadBquM5mNFvn/vzYbHV2Fz/S6/zKazsN7VhvvNc3Iw+YH75HIYcDMKTcVWLFopr
f7IYU7STH2B3QdiBgseXuNf+YdBckOIcW/2Z7nqlMFaQN2+KJzAtU83eMAENhg6mDipJi6Lg1pnr
cG3q+JbWGL2+CbbqDvCbdPtYXwjIJgOcGYFLiBRF5okAH802lgbCUPLwzKjps3/+6JIKdIlZojf7
kYkmoM1lK19LH7Tk8b+M7gEiwxoXnW4OWmtda1TZnIPB6lxmFTmbXCMV52fq5oMd1gJNJcKC3CnF
Iv8enni0nYbuHxFm2Vm5Zl+kYi5+wgPgUqpE682ZXJWpUniUb8mkOU3slam9jBSfzAxn299vvEvR
LtuQxoiUo9c8crCmJLJ/7X8NWq8eAeSCUvQxPNMIpJgJ6LfuOOa9Cyagazq6wQV+dE6MRy5KZz8b
t7KNu56sQfwuIlxN4lHproDWGsRAvj3KcIrXESE0bQqTTdZ1ryoltjzQgWakSvjxRDagUg30Ld8N
+r29UfD95aUn0Ym8hneO2CwHH0hHUg9cUcHutga4MOSbT4aDS6vtovz7ypDHlMXvrHHZDP7LjO8Z
JvEEJLrUiCxBRMPc3OCOPW4HXJVveoeTgh2MtZCfJA5J76B8iYX/y+grWhstfMk9lOIybscXYXKi
xARvG38WlB+WL/3/G35ZjGBmTBz/PTooGHuFO+zMZ20BhVLqAJ7VEJa/COhI0dKdGX2T878x59aF
LAXd/hK2LA4BGXBibqt7YA8wjCc4ARWbFjeR4Y/OWzKEz0QzCvldpf2ce6swpK3gN7DEjlErR3OZ
0WbDhFmfWy51nANxraEs1BW75dvP/oX6g6CKkPEN2d8DnGQXTKlXGX/Ue4mvJK7ZRGvSDNDI2WU4
bp9p9N6YjbvuMGeO9G9h3HqBDWW7Ppha3Klbx9cJSKZMR+wFiZ2Xh0QE9WaeweBuJ3j2fnWf0HPp
A+kDohrRUYVJeEWmIBjwJ/qj4glN6Mx0LUmaKPgOqJ+doKU322Z7fei4wuykjSbvIC1pI1odP4Re
l8Xx0AQotWeJL1RlFRWI0QoJEweMLgvQg/eIlEoJ+jj6YMDQs9eeOjbyY/5XVeN4jemCcPTmYJIO
ZOB9U3nm1DtoNXmUfmW80x/qcTKfbV2NmGtWIInPDZjhxmRcSHqCXw9jL5RJ4Eb3wzCdR9N97tvq
A2GIEP2K64S5cN0q6oP9yJP4OaEOjS8OHISRA9kduE4E+X/31b49pGsHAN33honKMiZyw7T2hLuQ
Tk2BGoH13jb2vRHr+amKxiJVGVH87Px+7Ifaidua9O4kYX5H1KIgJI67uuP2MbMXh8hgoV8biBcy
g8ooYo55iVF11YeRhfdxGtYUanIcDDE603zP/TYN0uXE+KGNBFDWEL6CvJyrX7OjTHCJ4BtOu6WU
jZSkf/8Jx2KXtvdIN5ilyab83vJn6KHTTVUrd4ZKQV+AKX2RVitDPSc0N3VKDEJ+GgQf9aaHPG0t
V0TTmrScHbB3PYrJaT23K4y6OZ0h2LIO7s4NSbSKkfU7oS/NnQzzsO/LL4mxAOkXsOObLcC8Ea/H
fB6GLzuOi27yn2Yd8PHSWC2f9Rav28kLSlLY3xDSD2A+XMzu6krNMyzcVK3+MBvojVOj52Arl9Oo
avZNo6cBMjZ7oNcSfRTZYxYeXwWg3YGnbjhQK0ZWG2IlKQhf5vCw/Ier/zHbou9Bs5RRkN3YQlnU
uSGnDGyCcrol8YrRqWBPJ1VrKxyTLr+xH5a/c/fLnsHWXmky08M9QBKzsAn9woYVyrL8lXqIOuY3
wUV/7vivA9t0coIXFrHn41vWgP0oD/r9mL0Fzt76frJ1kj59H1Ohik+AGm1kx6aRLGNgIgdKl1Q/
E3PnpdzWzKp/eV0I46kciVOKkKA3bzuTi4FFfzcQsHhz7yB4zUEmXFvDzeYGz+hBg1t9u7Rv+mtO
a1dl98VhCAY3l+i4gjtPTMQ5wZXcvEsbhuk6jcmzloOiS63rFoWCSkZ2EkeVatt3zOav1A7cIE4A
yKnKewRrJJEFYL5wbx8pUCKjRwD8K9JEbI6WAqNsDcH9nwkVdzyIXEB0cINyd3ZzTNoLn+JG6OQY
LeE2gVNbkJlRHfZMTkF0I7mFITYCHBom5NaH6OcC1D6pmooUqJf4g6SvsafNsRZtmdN6CTmm4C5k
OF/NxWSQ76sgD518P5fYB/cjYcDZT5zpLKn3uDEa4WehrXFfPhqmfRBV5mIXfHMBPYqpxNK/pZRE
cvdDtvqdW+oaXHa0dYTeMMvWqWsY6o6SsyHgAWG5eLfEVLM7U9FsvzH7Yy4i3xMN8tsH5OaJQcbz
pBvKUDLi2J2Sq0N9Ar9C0exdRuYp10iMATdKWA7lFwCiOrUFytWn6/opr8RvmBk2pygyH4SkZ1Cx
fhjlRdSCik6miIEhXZRMayPNd3zTqk8N8/sy2/WUlrxkTsIr3XLzqn09svvt6reUgcb7w6apoxL8
Wjfs103b0LYvX+4Yf99L5lHG7gg7Cz8egWdz3jrHCKGL7naqehvgeXSHekzt1l0MmMDxWOYny38g
3YzTp7cF77GyLJT1IYkwaLLCSUOxyO1Wr4HuS63bTfJF8rTK+M1Cqbqfze8X9JCMH9V6ZFD5v1S6
/eRtp5v5lkQkhLgnFkSgsGGAtSPZaLws/9g/Kfe1b7zwp5b/YQ8gop0x0bW6RQ5C42Ogd4QxSDn+
qeRQ2giIq90RKYinAPKWeJbtWkrUA0FLhlFc1g+bYzu9VyzpQK8ZW3rOTf3+OUX/frgyiYdzvq6K
SLTZ8WSvn8/y6rTYYPNFxRWOjJUBqiOl/TwD6Np1wpPgJ6lbEZuUSQEG77v2Xf8t32ipegIU/1et
M/rO9n4NRJ2QOLlHk7oAZ1UxzQn8wdus6TM5cU/Vb9eYeVkoK6sn/T3uWfVV/1wgMzq+BX1N4dI8
5ub7z0RWZNqc8JzKxs5FTm6hEO4ciK5ayivlSlduFlkXKAL9qUNDSwIi2tKQnRTSjP3jEFWZQAse
Ln7QgwsJz0hE+VDuzuZX2INWuae8hioMIgHNd7d4Q96E53TqwabzH86oxmrmhAcSYliPQE+zFpTj
5Hw36x3TP+i2rU9U6or25hcqygKCc25lqp3npa0Ksv10VH1NgjRZZuUSLFaaslpNiTT4y1KhGQcP
8MgNT2x0KGWO5VJfEpw2w7ZyKSMM6ev3t4F8t7kh734cDjAswyOxdC/CdYLnnjiaUwFGOwMITm2F
qOiYWCw1oD80YqSu0Y72vvUIi2yCzv0EpYDz8MrpYaSyphjr9IVK5bJye01zhxxkOKfFO+TGvp4h
CszM8IW3b7XymiMvK3fN00C27Qgq2vAxDZm361WTqavrjO955NgN998xR+ZAOWwkxwLJucffCEnf
5daQOEkoAF2IGMcBlyokoxh0zJUk3d19QyQciopIQVkfi44Rkw+Jg+9dcyDHuuZ3Sg+0opNPmzn0
YmmkINtronNOebZBAiWvKLJjHg9oZQzVFAP4H6y8/9de5CjoNeZc54DJOYqPaK9hiZ5j8WuGxJuC
ZNQgGM1PgyhM4kCFGpCvLAVcdtWMLT7KtXuw9uGTFTxeH7CjHR/ZuDqm8kulk3vEyEj+ZSZmF90M
WmS8XV5qOiScCYEaWwLAN9NjAnY8/d+b7ZSr1lUDMNt5QyaMSYZODKGILK//rELtWSTJu+4lKUWS
u1lVxdf6To6I4X0+x0WiiYrfZhDBIsr2qEU/W+n2TSNM+3I7Rl8jmisESC0aeo3tvqME6LRqok9I
X2pB2YmQAdsomXf/1jm2lnZyBK3uFJC8g4ixrGziCezi2XrCkyBbn3jkjjdmDlWrpvGJHjUJutWh
7AXNpyX5iPb3XDU6dRNLjbr8BsMab2yxIyhixvXA/QPpOzPHnEmsoI13J9E2GH6lTPKDUE4VW/LQ
OFhjicHKtSwzygErcG4Yc0ULgOs1enoIs2d5uVdp74BuOrIZ2hWASklbEd/oCQGyUMyKRbW6t5Yv
svg834v5fEkYnfxx5C/uvOF+3gXtBxxDjH9reFx8RqqSwSpiVEOjoAHbaXIPAr9hzZOoxH8VKpt6
OQ+jDBXWIIbBl4H/83T3nmAFbyGqfwcam0A7sac0KNx85yc/VNCuZw4koaLdm7TzHaUm07SHilaG
jYEznG7OD4cAPayw/aktEdqFVBvDfX6UuB/5jxJ3mGQoGDsyRyrMnB6M4+6Zlki6EiM5/66ApCPa
9iF4uxQXfVIAXiEzqiE8LYi2Vixp5Wr/8hn3yLClmVbnxLuH3qyGBZ90+CkB4aYnwX/yXLR/Ve0G
fQLXU8Vs/mFEK/bN+l0tjjhovIQFdyj+kxEoxgP7HeVVFdNtWhps1zVOnky9InTXkkk77c17JENu
WDeSvU0aixAZE3quYxGEIqP3Tod+iKHaVaWEpkANTAiKBgbr7shS6oJ9JnOza0mEBXFBPFBb6bLp
FZK33ExOkqAXC09+PpAU2apGrWjuSoQfdYbYgJnqUI2FDWppuFKFFYcXCBOqhbH35Gmgxu7XJqf8
4zbbYq/TLmD8KaXWXPCTT+wnvZ4r4mSsRoaYt5xdyTvCuNppJLEqjqnTz1cLJfnUIMoQmOdMc1XO
bp0/jZHP7PxvMFeE8MUvWXPy3RMTIJG8QLlkXvLgGxaeLePe1i0WHUGXft+Hn4/XK6RGzyYclXgw
3ZaH6jUDJip0TPtBpasHDiKykEaMefCPpqilci6KI6bGCQH64lLTsv4FioBvpkNh0jEN3WDaHJ75
OtTIjnxHAycOSEDkODxK5ftwgd9U+7AF+SDtXFCRwKwUjHi9v8/SQC/rrakjVDZy0UvmZgBbqemq
hf3viWb4+hF/SrZTVZSES0QCPNSrtsvjDJDC+ffo5o8tyA+tFxutwCtKa6RZjAtCPNs64IGR/b9H
VxwoX2WlKJHH4IrXhZjCyLD6s2rm7iGhoaIXSqfbY0jgwX65B56xviObCar/NpylIL+NSgELUiG1
F1vsH6ok6CxTXtYKUa6KDHnOD/V16upDiAZFob59btv+rl2wKqSF1lpX43VwUEEwlBiVdQUWcyuB
PTOxt0k5tx9abcRt8sthtRUnaOzvMjRDDi42xsqtWrwe48Pe6LPcNJsouB+xZeaei3cIUUFk0NAZ
QwYkuqmwi/jILQTWQbNs3qN4vOzigWC/1sXH5we4Vff53Qveba17Rfuk7w5ZgzBiBaqSxuITOUZe
8WizoRGBIvoaMnRcI3pjD04WGeHF2JFwpGNDq6/TNQZiIQoP8/BCJPURq/Ii8DmpSCZ3TUxwdwfR
PyT0ffIFykwRwoMtR8BGV31/w5nSoSzRT0V6mrGBEXzyZ5bemKZC9VBhgeiqnsKXTj9whiyEarDX
m3kt7LuYrv/p0g4RVF2+oqm/diHekExVXuy+nJ1LH1SYXqr3gK94s4BYBxeYBDmR0LnmD/50kiNy
lzInraCssKcWXUzoa/lvqW1sTk52iDTYBNoe17Y/mT3fw9IQoVMpsjJiV3V0Q10JQQkFnr+5qKrF
4Msx8TRN+2EPJZKX52DbNWo8ZYhDWWIU9vEiyKkHBsUyIYUqgE5zhBlHzWaZ0MJ3hII5+Vf9evUd
02it8m+9MvJKh7I0tcD8m7rWI8TQ2ityiWOiJZNISxqH6J5zrNstA7ZEluTkaqqmHQX663AMDM+M
DYxQzfj2QGTscmP6Ih2uUAUK9Z30oHD20gK7V4zhi6QMhcHjrcc05K2qvd4hdgiNCAyFHibgXsXM
X6snLy8cwKKr1t9VgF2M4jIAvV3o0TZG7EBdXYdKVMwFB89O3lkClGS8qWBmKZxGzwPjyHcThm31
Vwgh1GLEi2HUkC0UPPGGZYlAzAT/iUCV7Bgzi2R+QBgX1tOegoT6I61wqYeDRLRjjQ4UDyNvJigU
iMPOzG9Y6fyHkLXYuenut/ZwNTAKxws5IzlAg3R0XcorN3YpBtDCgjFdkPDpu28j4OAUxLQDae15
O2r0I976QxbTYW0jTAbZOCdyV5PoWhRr3M4e0jL3oSG0LJQOHEoFlAafpnoDW+kZ2utcjFFEjcG5
JxJ8wB3kT9Rih3phAqh9Ej9mszwp6sSW7aPCNawDH9eeqsFCtCFMiZyINk8f8W7SeMCPnKBXKP0l
D/V8c9Wj+LwWGJYWGLJsb/xEowe/Hjx1Vxw2XMNQ5b0x7k4r1WTGVrYae4RkOr4DzGAUeEVoSUXo
2ftcSJYwrgJA7JfGUaNWtIyC2ArWRzYNYGpWtBywOQ8PPi/iUW/x+lrocGNI+SblssRX7ou54U3A
Ye84GOGlkKy/ZGUwn07jSYu2T1nKCtnR+LSUF8zSb+jnTFI3931MdfZMNBFoVCfL3eYUwEIJNps0
fKNsxu5w18gJEuLCyNKCCo32/4r9ms/m1srUDuFIPliPpO4AFgGEFXsQdFLbedfBA1Rb5nlNn1ma
FApP281JW2HsJvp/uL/FATB3vAu8cPmLKJyy4fXpVvL5whh6DpB96NU/s05nUZ/J+g+oYAkZXOeY
RdmwvkkjlD7JSSv5YG6X8XYFFVohAAqyrETVWJNi71jYgTOOu2d4Q0wOh0CO0LGl+JAMmebG2nvw
xrAkPh8dEJpsirybc+4xRzYwuni3hB1iv0FyEMln78YqgpbyUeVOOQA7EgVy7Vq+XIB1LtVIATis
MRBwXejbctlthF5qG06Oa15jb/MBwuMvWyVmaPfoGCcNaPLLEy6evGLri2iEwIjya5dzs4D/8L2F
LCf3LOzHoGKGB45j0GSGldwLs3JXLoKLwEiPjgP5dVnal56HTrsvE77XUnaEihXEddprtwVCIhfu
BK069jGDF0hUr9WhRK8SaR7zigok5XE8fnqs2Q/SIqn7Ui739geogxXwSR80O4rrq9cwJfvjrt5R
O2fU128LqUy3n5ZtZNMSf4n9nsTFdE7Wq1qKaTVdDZ7gDsQ8K6uTfTyK9A/aw3pc5oaigyS0LFYn
bzTLRQ8VaPnCCZVLdUZ33v2FP/T/0ljtGA26d39Q/gYDc+vGnG/QEOq02j7CvPi4S0FqpGVHc7LA
FgCPw1wl+85mINTbN45KEGeEV1hVdHsIDoS4Z9iaVmFfE8G4SVAemqOhx3/cvQsXtLU2rKHa8ViX
kmGQY44Bs4T/NYzq1U3cbtRi6CASoYl3f85zzZHa2cLgtAfMH6felxHfnVM3574WdWSFizQaJFoo
03SvMC/plpQhtd/VvJDFl0ntwYLBNHUchlVIt+DWb5wwitdMfi6rLdRHmO4LtbHv72RE6/L0qZFm
CEs+NC8TToGHK+WkvbzT+dymwvgVrh9mpg+qArB78ikt3cW+ZjgQO3/cnz3hfJJ2fdE0wLwB5j6R
Wd6qzBRWosOsgzwg6caJJGrkkJh8kojgRhE9zgkXxEMOH20s1DKHQycXNMxsvjolbyflPpASsG+7
R4yGQmNK9a+6EWs2TWZcc0vr9gm4nEiIMAkShH4luHS4v64XU2RsyPm82p4dHi/YFfnEfQcS5icN
AXjppknCzfO47TH7c9Pn8+iUe+vEJQVsXqoywhM72RASCs8bQCUTQ1dhIDEVW6eoICEbisVBdXGt
BFrUbs0v9PhUdAVO9OGlTtHJvRKknq6ZUcLCDV1DsCtUO3BiV+1CGYnLC4z7TcHA/RUr2WO5J1Zh
S1EBIkLKx19bcJYRduvxC2gNQR8Tzt04yyqOeEHnzKiuMK58w5iSaYIgX6Ua5s+KVXpst1I1ozPM
msQw8lTsd6DBdYfaeBXJsgkYAXg2BOcCIuEncPILNCrTsOyXvh9ZGZFigvLN3NkGVQ5ba1eDIYUh
ZkXl+VC/MPNqIXV5YcfBSEdSxU0Hdc5Ket7HruG7sdKUk/LwGeR90AYhNIacbSNdOBFjF0yRVeLS
C0SJA5ZHFGa2SNdxPskKvPz8wiQgI6aDnPcbdw+tjyNtkQ7GAb0PiURD3CxTP7S9nwXo2p9sNhFs
yJCFcNqxf9lrM3ft5yBK5o/LKRXqDF2zQD9/kZa+xqamxWaS2SRKFD356cFzntom5fmkrd8rgKbo
SL/3E92iQKMz953UJLcOqPPwdjicTF9fHohJarPjMBOWUOi67//6iSCWISawJEOcCbG7q0Z+doab
0g/i9t4Z9XwiQUQ7vlrwT4t3oXbUafUymY+hfEQkLSy/wF4FAOf6mLWlAtRvXI7OyGH6B+/BIIuK
Pkav2IifoOw/VdXoI9+vsVL9aayL2W/N0Gf7SQtjY3cQH9BW6nRSuE0T8WJFz3mEazAw76FgGqVI
R0zhUIgTsU2omCeUH5DpRqkoEB2vX8iMjhShXQSyv4YSRJrM70zkfOSJvCI7IUQLe/DM4EqeVMZd
QjdLZskSqdR1oILEOd3wXnLyzrztSlxLOvv1mSZMZqcl2KP3xG4MXzpD16ip6b59zrvMd6KULVFT
M3WJX8KdZo2wKnRoECXM6iDpHuixAMXr9+8w+F1LrSNNsIiF3yPuy5bThO0EvrDUIONcY1YEkgzS
4DVwa4qb/RwEKCNxly1Ldj+SoVFO8g+OV//kH7GGguJjvNm99lT0xvvDkBWd9Aq0hlTRqpWLky2s
njBlxqDk7C7ikvu0negD/1XugA6BQb98tNsLBVGHxluqdd+EeagNkszcSLWPy5ZViUddYBCgMCUd
B31a3eb0pdlQRnpzcq1LVCE0TA+R5PJqNrrG5KR/TkSMFH9ZxLe4FdB4+tR7z2AATUL/rCF85Ebv
u/Hq3Ha6IcJwct7Jgpu4AqTIE3aQEJFSClj1OeLjLSFWLDN3+TBmZLcXbq6BOMtVBQ/MhWlzc6jb
52xWuxQjsXTRF5FfRME1XLfuAGKye+q2jah6Lp9nK3P+1/tpGPB56p1+RoDQf9ER8aAdfw2WvXwa
mueiDfvdKvaE7zc/TEMssBxhBUKir8lEEk+IY4bzdDwMc4YDmuBNi5BkFNwVKr2sFQKJLZ4Nwf9d
SftLxxvVLZqXPdZ0JLxxF/KGCsUrR5VYBV2Z0GlQjJ3cnE3T1J3UaG42gCpufcehqXIIXxmREYVu
ig9O/TOHzipSqHcnJrzlY4whID3WqsbEIBFx7tA3im4kWRMwk0Vh4kh4pfnMEUGa8AAkWzYxwjx0
iytTs95Vx8rn5g05iClb8jd+NdTqslcA3agmj+ahhNw8nmyJm4e9N+wGmcwJe6kJ0AH97IymbYwU
fuUAvFO70gBErzU1WNoWZ22A4VF0OTwhXSKb9/lN1o6orI/tuBLe43jkBI/Saz0i85F4Raks2wDS
/oDAwhFnakDyDr0jbkaLbRkFgGr0p79YlRwy2TQV8Moc4HVpOUK99OsELRKOb/mbeCYBd1O6PrKl
Ij/dSihtATRWKM5r+Z6O9eELAy1tLskPhLd0Hz/jfD7mBEFbVydMdOIK6fPHwmJN+/UJbSb3J924
BqqY0icf9Ug3YibdgzL93QCD+uyrO7AGWwM9xkFXmtS/pT88bAbwobekfz6QjuCVzrNTtQTyr6to
kAwdRMt1R+IvTCL9hoInzjBStXVBgx81XXwNVg4MTSOfgL0HAkZnp/TRJ5TNNqmuIlC/VVt67P74
vGBmS568MD7gkyZUUAiL2/L1LSOjgeb7G1rhFV8obpyVt/W4XzEBT1S79EaBylU1hKldbTBQurB8
rWtCVpuTltuje4eW4By+jpHXVk8ZubhA326zCJxaRAv7ogOLH/CBiOgSgFDPTJJec/0YFxyfqP72
x0lcYbxAY1CW7aSTEqo5KgmavAnKuvXeFA5Pk8vpWQ6CyFJgt7HHl7agDpGcfMhMoomMmuwoRmYH
Pl4iOIBnPufkHAfdcdsL/uLmW21dpF7qqS4tnh75z7WQljlKEoUl6xwCy8LO1J4Ku0/JfFlWVZiw
x1mmPAg1Ia95WIE4nZ6H2RdrAweZFupbPJmHjOh6qh7ixc4WlpjC0qr5rEp2F+uRdh291aO2iMUt
Ifqw6vZQSn4dIOgvyt1SpYKt3GCzVHw0XBv16UfaF8Ios7ZqAsnjl/2NpYTvII2IkNsrv5OC7b4C
YlOWqATzCQ3BOshUEpX14gK1nnHWIgrYgwSi344He/dFrFHYpo8MuZhWqvuZneqdV2tVx6o/v7gL
LpB1vFrYoX8Kptn7uErfXm2uSSlVR31wyX2RpC2pbM60gjT3SiuGrHaVvNJO9z57lzOJCtZoN+AJ
7VmsGydv5FMBEUijAstE5TgpCVEXXBYwQh7KIjbUooMgoFhGMGC/4MFMoQ/H+QnZTUTjvstZ+PwL
VPnQ8oGhSWjiElxZkVx9wpSazRgc5l5Mukfc3nl5vz0hhdAd8Vsq23/3Bg28I5WiN7eM0pZTrkYu
0hKd+o0VBAFf37PnYVTdwqb+7owRFuVIDvxr+nEGFR0pYRzPvUSvjhhf2clwK2d1gxHrCrZPjPHu
hMNCdVxt7S9w/LielU29Jc4bUVI619g+LAjTT9+k1rximiNN5rb+YhEs7OycpDj76oNgOE/qCa8I
+L4hqitYZqtEpr2MMH809gR+pd5f9wlcrS0vcgZ2xqCmBUMK64p9GvLsTcIiHhl3IP78//DKDyQw
UsvW3eqk3pvqx0O9ycRUp3pWSFA69V+MtJ3DLTO24tN3VEq9FqgpmvNJSYlqfRkCdUE28XmSsyWZ
6rD2oEmNxqg7v/eODZZ2qWovWc7iSzR0sbw6Jrfp2QB3iOqNdYs+1F1Vl85qxWH+I1zn5yiCzKst
wlwUKpmfz+ORdkAAEH9i+YbwplPQoAaFR5G+OD1AA0crvAC4svbKjbfcu5NyJTYMQSjUGE3X9XPF
MjFVsNQM/u3uqvdhQ/ciX3pKNRAKGpE3XLiEXGK2XZU7MPGzM1h9/e9yeWw7OvgKGJDcWNFdx6Tr
bSyYX22VxwoNseU+KagK5AKV1et+CATwzwSMRH5arbP3/vGxV+J0BTBcehgvJMNgAvlph+hWGQ0Z
bkzm9nSaZ/ykFxgRxIT5pFv0OO3azIJvMq0/ha9mrJRseke06NqVN4MTncvTbnBEvGNDkYiyhCky
LdPbnnQ+1HShfoeLM9Ni1kYeY6hAfkANSach1WJJ0N9ZD4Q/VkUlkQ6/YmAFiUqrTx6bTU+okV+p
6H4Z4Mjnz0JJkCivaArfWzwZulb8nRwiQnnErc/ZDsSPxGGNEKd+fC6H/hCY8u5zcChSDWeFOVlL
h8a7/Zw8PQ5xwYDr0l21Qs+dKKP8ausRUrlSXivNQ89bhXH8wiJBZNinnMShUQnocuvb83rPmTW2
9DwaEW+8zdnEkilhMB6G6dnyFxthNFb+N/gLDvghYapBCPsZewOEp7GfBt7GNmRUVbZYKVOOPapZ
hqDsPMdiWhaOIo/+IDF2My263nS3/bRmX3h1SZ10rWLcKKbJkqGHFglK+TZm2CllKAJ2Au6JmhcW
VPK2UidWWzQhYhcpDJQv/idARMySUYSuqz89dbNcw8ZINMcRuv4Trm/pNni2K3W7Bvacx7Z+NVt3
YtV04SIEW/pLUUvqApedzKYnjmdMB7p8jzVCESjQWOMWTOmyZR17eTwD8NgSuYFK91cDKLGKRMC7
6vAJi0xJm6vCLc+yRbcS/ahdiXuFjDqtZ6wTtH0T5OPqhKbpzZj3x9bELLMPYmpqPIDiWaOvvplA
P1GMQ/WT9kBnPVVKVQ4FAjyengTuEk7Ql4cDMV1Oa5VBBajgLeTa3bVskC0y3Zbw8CGqE1ZO0vHI
4LZ9JxWK7nAZb4nRq8QH2KfwJWnocByupOsZmkXPMHbBKJlfc+IUIva/qSzSJP2HfjJHhRHtK7oT
jzvjjFaqbL616EkSVFXZhW7SGrPW8bcPMgNGwkRzLJDW/xpiaweteHfYx6O6j8ctBtj64ZqGrkb/
J6YR5fzJUiYC6D8kx0gRgPdd8MP3R4dmXMRWlc+7essDCyKnlBXp/xPrxQQXoDtvOgj1ZPj3Yi1q
s7WTNjmdu22V2PBgzz+u5CW/6+GyT/uoxHhP/xmKXPkIq9UkFQNbFn66/kag+eCxgxEOnvYKmV0T
LIz0f7vE8EmPeacAU5stq/4pCWlvycPRbApurF7vpa2gKU2A3Hzzjkg+kuwhfgTFkk9kde92244H
DaXt7PGp7hSmPewVmOL5Fy7tQrUaxsTGfA8yj8P/RAHdRtYIBDItmqANcWGREpl1haSoNnH6ZAd7
aL334gPjTq6rdgJ9KRv7gelABRujBSC5DSGSbMRs7awqrbUhS0Xhcd7KhvzpcFNnQm9WvzavG0hO
mIfCpbLZTb5Vi+LP09c21A0qRKwDd6yLmalRAgxV2R3LE1eWkcUbL4tbZZzjiR7nP+FOde5Mcd7M
xZvUMvRONsBeE0zahZGTrNecKZe7gTvYRjpXFjTN+qkmDZ0cuMpVIxEBI/c6SavUoEsLDzMml7D7
iK4cJLIFcRYneYkM1ygcL/+23jO7DbHqQK9P9eByvoHqvtifsqjDltILxXASkcls3XBXACPKBy9W
j+jEqgT7QUrawUi4bCyJhD/v+lgUvc4k6aj23QmeU7diU5DTWTk/9R/d7CjwM5TcYZ87C+/fSpHV
gL2vMXz6ZoWU9N0zXCENQs1RLjkzbapiLCIfTdElnKRmjsGFjWYZq8r9XjdjGLfv9ThBbTY25U+j
TSEQG9VYc7VHNQm+wL2RmU2EsCHkMisiJka1x/x9dJqZKizrAQSvw0K9FmLDz72tYJaIV9/PVvwJ
84tA3X9Gqogid/TnxBGpsXLMX3mjboCRT2xMcdtL8Gi5neTYR1ZaKuLUJ2LLq9JbieNUE67HZueF
+cSRXJI95k+H74VCT+KZ4M3txPsqHilqF4eNNsjgR+b5E+RE1ln02UpZC4D36341pUle0JgceO7T
JLv1wWlbrepeV9d18hvskuT1ojp75WShR6esD/ZAkDDjW6MTIroSDgMaN1mLfWXfEv55L/u42b1O
fjOw4XaCX1ez/ie7zt0zfsb+TC2PGbbsJDpqZQNoDgm+0s/n87S/8RbVA9QLIbUWiJ2QXUYHmnNX
zR+1viD61r3Yzy8QdPjgjJ6EN3r1W7GHdkcn+KISuQsVkrvv1R7vC89yFa9hBByMJZN3tvplMp65
x1GknbvUaYWltRF+lUh0z7XJ+utWdQll4e3XlPD0iIHxTAxvK51T5bMC3zupfYwGZ24sDm5VHhDO
ks7Oa4EWqhX3eHfG7GeQwe1ulHFpUnoyty4uKncw++F1MsiNI9UMT3Y82gIBxeYEQAmWOcPkBAX3
6HHg14oaLBhBbUlic3EQaJ8+ERVpFxSSX4f7Y+89SiPvFveACfnySKW9jHbe5f3fK7MCJLUAmGiv
gt+Lvsxw/8nkK05AUM3S77XNSAmq4OI6GCJzf7pIKI3WZDQOvnR8x+fNtFhVb3VcnpL+M+hXeFxv
iPCqFG1Q14BSK0bXMS4D3QM5/FK4zHMDPUSnSzcGf0y44yBBao8u84PVCC6/ajxRj+VFGox7/AGI
VxLk6x74lJJc8gCagl7rPJJStag0tT54NhldFg5IjKtDX8byuLlrV1dGRJgW0copEx6FusNambMr
w/AaFbbg1chBbu8QsGC2aigmGfDJspOzo1PPci1Fk2vgkgS2+FvUnbwfLJEYyCBPCHBCqfk3HPXP
PXFeCnR9OznW8vYapt5RvwEQt7xC0QDCNSis/9NU1Mx6uRsHdg9O/okEKd1fAiqaYzUM1wb5O3AC
fcAze1stR4BtFh2WF5esABe3ZS8Bxd2RPc4G5FVO52JaOPwSKvx0UviWn4ofwF+ctWVlGxUjzQLt
SASybMIWeuTKdWz2mPnWA/23BNklgENToE/UaLdBtprn0suICzFtswNOHx2cCzmPy+yJjgI2KWp9
etfhnoUbC/1bIDEoHZwG23HbTNj6/rhMPBayzt38XK07uHc0p6ZEts56T2Xfu2TcRK5nMubgREwA
nHlw4HYsyK51XGCX1x4PM1URcH6IXwi/bp5TeXGtDBdYLNJXoM+BHfNgvtWeo0R3M6WVKaLgiYsc
IIgqytBgeme0lSPfftKTVuuII1yHqzq0/Am1lisR/pRBiQs+AV3v04QXebsDVK0yD4Dl7V5m+2n1
riMB9aKrAfEy8FvgOM//Wd1QoHF4cq3K2LVXnepJx3XYXyzuuqYQ3TbvKpDqhvSLGGvvGI4A4D/a
XNBTOzycBTHUyFxYXdgGfOQaOXqH4FEQaCF7bz1TV5BD9Mndb5au4GTq9z5cQ4M7M35ms5sPZoSb
j10ViUnJmCExU19y5m7NH2KBCkHiYkC3KIuckGw+tDYXTCx8MVquq+M2Wemdb6B48J2yd/FrpZri
X3f7oi9yjqGR2Esiqxw4sz6T5aYDO6bqGvRgu0FhWYxPx7yuBRLN2J+eVUPe1AQc6EUXZLDtmIu+
zb+r+rfVE1XEPRyuc/RUrepL/3ZRGTu+9a5Fiao+xxTMG9FwAOaaSztO1wlHLClup6eCAFV058j5
UhAwOtcn5Joen108Khgqiv8Ab4AdSQ1mdzGEs0CJ230eklI8vrmW9cXKQLidEwDfVLeAkTcGNjbT
VMx69D+Ejk5uUUfABynk751u4REZXdOe2c2knA6uEJfuMryEqUb9pBXt/fDtWhIapFEG1JUpGdc7
71AFUoDRQiqLucaJKfpwhPp0tmJm9YgIzg30XcJe2tgTT1WAqmgj8RHoYL/FSz0UU9OfzjKCI0Mi
F3f6sp6fFQ9mSBQz9tA8lDNrSdaWR27aiCL+jVJ8ebJdthG3MP5vdLrAYsBtMJYH4kfUw3EJk0Mh
VENJ8x4DPyKuQxlJrRu/gt+2mnTUERKZbNF+RAad0lX2uTm8iQZZ8VF3oRZKUdE3hwYdWtDkzrKV
M0CcPYkIokwDqf5VQAqeI+GuflRWis1t6kadMpv2g9BB6itMUXjxs4E8mQtNvjZqCJ5bh6OK0ZEE
H8btQVJw1GzNJdI3G245uwgbHOyO1l0U37K4EIJtHcq8lv2bzgojTzUmvE+wmkon23/bo/VvJGeE
wsL8VJEafxBMw7f3z+LR4Tp4RocNw8FoD4K2FFo4ptjbNS7UIVAoML5eSTMvvcxyEDOvY9rtn0+Z
uq55rN2uTAzghhnw8ywNxezcMfA2vGeyZdkCg+s3eWrpgF8X+Pq7+9Q4/57PegePmtj/4du4DweO
h+T/6mGfWlHojVs9MA7stxk+4BQPQthSLyzngUE2uJJf6q+fOPRGWRYLe4hIAte5VA3+Xh1d6vGl
x3fa/eC2eZFb+safkeKb8fpBM8ryF/GkM+G+Qv9mxVHKv3LD1gB7RL6ihb/4bKaAzu0Mlmk5exJU
klcxxMrXWVwJjSIkNHRS8axg3aH+sMq1bIxgHPkZWRg24vTYNOnaMOBWhVUyP2jYu35F7gsvePA3
Ayp6V+OlFRE6MC8qBdikHcn8KWs0kPyg1qLLRPUjx2agx1zLAloHCQQ29uMH618rrkkEKRBI7lGE
c2YGjVlpkbX0QEJn/++JuWfjMqLjVUyc7uVziKTv49LRnNuy3fkUzO6QBCCWFvlSl2C3Ads8xwrO
fCOvwNoqXr8Drpe0ug060u6WT0EESkWxn/8Q6GZkldfBHXkiYUsd3i7aUk7xRPY5I0n5vlrd8/do
WSsjP2Rw2QOOvor/AzDfVK/t72g95Xd65xLcalK5PqNBgkKzSJZY+DO2QbZjUS5CYwcJTa5rSMT3
q6+q7wCA5RRkVuH0TgI+3YPe7A3JGrr7pTS6rQJs0D5ulw1yQGKzPUeBDlYNht7hEZ1rEfXAj3lR
yIK0thdUWWrcBdy8laG/qNi7xGXNWCgdg9Mx2IdG3weGK/mKy6M9Rw53ufPB46eIvDe4cFEBl6gj
0rzxWZ7B13rJQLu9mhuvloulftYuHhAauzSL+HDz6xChbJPXklbHrHz33cQRFoW/umPOJRFdl+i3
ibFwNyMRNU9qZJ5snUHihlQJjtiUaGr26xlyUCeh9aj0j6arq/SdkZ8jxw7lEACuzt5mS31WDMoe
LUWsO54n1XiXptaL113pmlyHjpqfg0r82ozwA7aGM/1Ax11Htl8IL2bi9jFAPiUW3Rgjxv0m8yUt
1cTynok1hJKXfc46xz5JdYyzZTkLpSyEBsWEcnYi5PhV+CqL9hPQLNjvCCUz48BJltUDEGmH6Jty
KtlK/rBfW0COR73fGfmLqr9DMuIfU/+7nMSW2nDclug6kkxpr6CajmHIoBgi7U46K8oYzZX2Bky0
JC06Jsmo1mUn1fJ4A7R/9UYhnH30QYF5Op2NrTzc9TuQX91rQ56EarGuL7atIFqtzMKbRFQFnSW0
Pd104lubg6ClnFKW7PWhZosldUChxOH10WqMkyjwm257m2kyUSaLyjiyZ7MvUN8V5gbOD3cpxEen
URK+Okm3rtR32qj+mhmBYf7LpaDnp8yp9KYJUQ2XqhaNzkULINcPhdN3tm8TaM10A6jVow+SqHOd
roPlMQ1nDUQQDw57cFW807v9H+7E3vmN1Uw52333pLJLmsLlgV0FtDQi2PB3LBwztoHM5NXPAffI
vsJXU11ZKNxNqhUw6gcyk7E9ZtuSFvHzsYqruGV3nm0p94u1OPLA0HYcQG5Wf0Cb/hYJ+44swfQv
i0joNdT6gjPobDHmYcKmE7P6qe62aSAn8CeZVOfsTOnsjFY0z6argKYJLMiWp87Yq5AO+a3+pPO5
YUrUk1Pzs5KBaFwRJ5SXs1ZZbGCh9Weoy9n4f/MljUzUNCWCYIimOjUTuiXFS2tX61bUzglbv+YL
scBxfBx6efYcSnR3pMx72sNptrA/KO/7JhbXsPLduagENTB7ttm9m0NYOUFA2Dci7nl+o1jaaQJ9
cbWgpoB1WRrwXzTlsec3yGsoaOXUt3nJDUE3wtu1qCd+E1IfYM92AgsNj9Q7Lur+N8uM57KfeA6S
Um6I+i8ZdAHkRAfx4vJcpvlf2PoDN3lIjzhBx/mfWYSl7likxPA6NI+isqT19nph+FCgR6Gs8Wgq
8+RFk48bdNQfFq2A0TryxJUs5UXTIbCfHd4YwWr1rbFAGNdTxqmreK5Q5V3MT8No/2gHS+w+bJcN
jkNvJk8ZQu7V677waqU7dijDYyXzkp3oXLPCdzWkOI3tXSxFxyDGTCiZPlS/HFwT7NTxI6EIsOdz
gRmAVuNAAY8ckh1iPLMOIDwiaUc9L8P6dWySLJK0TDF3EdU3z+DRgHjIziOIFhZsKYqqwjdGPU+a
8d4tBHS64GImLH85lu5pNXm+axMiJIXmZx08vYiNH1VkpgJw//QtyHghJfgftyg6F6S4PtGcsllI
QcfhZNZqf/zISvu4JITRvMPxJRea0/n6KWawRHnpl4/10M3mQOCJUr17SVd2DBZlJo7lEwFM7kvx
KV0TsIdlQzha3lqiTYDecIcFmT42h0K/v5sH0s3R4RbCg7gRMfdzj0HEOOLeDkn+ORCjLxRc8JAF
vrYS4eWvIeSTiD58MYtgtls5aP+NzllISY1R9+seLH7Zxq/xaMAXM3mn5lJi5sn2A7IRpg8mgFMK
s6tAzqI09V7liISImJxx729LDvdTQYC0RK1nrkEyyqjj1fJ3pMgb3sljIGMtQmDsSzOCrnAUBJ1l
/fJUTS84O03h1TN0VHdSWYiahlulXjmz+eIF9+v90LLnxNsVaPaLCjFnSoe2K3MblI/WSV6PzjK9
n2QxNiJmgl0/AvBZXfiq/x6VHveBIy8X9M9g67ACOVzoFnx4ZAJFD19GRq/8DGSm19uThT9QVg4D
CqQHOSFgP7dd9jIqGllnW9MhsqYr6OVyhd1w7Yt8guZf00WR9aooHSOqAPtJaPtuESvXmaY6TcLl
jMoz5mk6DjVClbLth3gnbG9YJcHJ4RPnMrbcFoiLFdxgSrFpqqij4FwCMpYqkrlA1DM/yiImbEl3
p9xNnZ/2OcRK53dSG+Nozs4uN8P4zDJjXh8bVIZccO4RsDqiTKD453l8LMYiA83LnO/an/NBWt2X
gzk4TpQIFpu2GlTafLx76CnSGu8FVIVVx0h++Zt8E9JP50Ho+ZxQrSbbeOFixMR1rWvaHSS1Fpm8
5853UaHcSORtRrw51V0nYFGyfg3qzektRhAS5GU7MYjtiqgShDemnNRlXLwpKCCRMIdPP+f4zHu+
TLYGjBC6HN5yiQ7pBoYLNsR6NcWxbnvxdmp9569My4HlS56RqgICO4CPEAZixadeniHoseshqxeI
LzoYuTHIlmeiKADyKsw3DQyb/9O/xThStvU/jopsjjKvM6biZQ0zMhmv8+Qu17zKQUMpzESWWcuc
U6k77lrelSylr0pYM9GjULGY2Rmg7BvFAEC3viQzrgG436CyhHPKmElb5SpDeOFsp9J+ujgPGTFM
I3QR+1Vdhsc7/aowWYt74jtu7G5Fz2u/fjzXnqy9PSFZaC46n/CTEIgaHp121arFd/iOeP1+qpZg
yXmJnlwZl/5cmAttYtK+zIKf2QSs9r45PDBBgyhVBViRjUQuyMmnX+rxFe7TpZKj8t79aVIUK1Ix
DQSVMVc5lUlbL87Iw+UO5Qoov2lJ0NzSB/Y/0zHeWqcVLYJ9mekzUKMSWE50gm84f+nzPS3MzayN
DhplxnKMEbMbJvmYbC9P1oXW/KRxn7D6xZY3joXs1NycOnablld3tMX+wrcDS/5baF9nAH3p8P6j
tqEq/muqfl/+nx0pdm522SXxRUHrWWO4jrL8DEffFr08iIm/jivjnk5A4mE7j1j16FEQEhOKLv3K
qrWe9kvtULVkbO4e+Xr1WUi7Oq9zNH1oEdqd+QJM0owd5hQLUTEzAd8g1SJQIqgey9r2VFLmkO3h
pzMWDCoaWf2ZILgM3gra+ddmey2+t3JM5H5z0L9n9MFJ/34mbtwqNlWjrX9GCdcBHdnJzif7Z5di
7x4l2MHtyp84QU+TYpy9fCkxRPmnWUUZMWtvzo+CtnkvdptzC18zFRmuRf6XmEcZHray6U9Km7KE
30v9j/fNvKKXMgWKqcIfg2Wqzn3V1YTby54hmuCr0b6uZLg02BlerIX7EeV3cM20xf8tbXsHfPyc
JRieU3gxBtfVlciY+5EepE7cgw2MT4XLWuJ6cgYlWvZYmRpl0a9LF9Y1BqyGlBUzlvUtOpHe8KdX
n4pFyxIv6BDNFge+8A1tz9V31pfnSboHoLIBnaviC6CGkOosjoJzt1rvAn0d9+S2b8IQWf7k/cWg
nIqSTpTZH/Boa7bs5mX1CnZwRZZrlVUOqoIDAOIkQIz2CMxfWoYo+/TuNLV6/tIWBUuJj+SxuXwz
fO1viv1HnRzLXl4kGOLfvM8mNPC0xJ+HniBLHIBu5vCCSXPb23mHxrm0HGr4srWDxd6rJxQjg1oF
+XXQyThvgaBPDnZBclyCuEAC0WQNRdzGVepA0TK5cgO9EGTw1pQ3X4ahoLeRX6TGPWgOB7+hRN3R
GK/9xtNIT0HeOqYIvfYbZiLq3gn135a7HjsuhSSPSKGl+Nftpy57KGflNieDDLkESfUClAVA5DmW
JUHzCJxeZ1BpFc00QX0n2cIUeX+SkKHJ6OpEvQHwHPx9jrUcTFPkPK6ugR2yKAtdMnKTr8OS3bFi
4r5TRkf6yMsONeKx/oJwWI2s9T0V+up3tsEtCCW8636g7O8CaGI5cVoUjB0ljhF7S5DpYM0W+SO4
VKbGvT3b8WxWXqFgkU3YHMRVXglCkCarznli2/aI8erzUAxE9i5e39wSZAlelu5jocp29zyJcPZW
vcPP+jfXublF2jMau6/gljQICiFNxCxfkgnBAeR5lqF76e7+k6xNMhZ7Ke32WvorcvhocoY1m4db
DHTqPQ+gr3GLeq/MbUoRpVUIiOKa1IbDjLi1dHTqTjSUTWbw08AXvTZ1GRP4QyRtok/x7lGJ90VE
I8ITejvhaLq7kcP5zALNOkFQ/qzAJVM7WPitZHJpdTLDJKCMjJwjILz2opdYvD+ryVf5Un29Gpwo
ujQUBoa9OCb4fOUrYJd4yyoV8uQ2MHo0mDQX9RJ2S6+E/axbdwPEYmaGtTvwyir9YcMkj1LJ3QPh
wQoRtWOj2nEANN11Te7QAhbRyRuEvVXIF2CsE81EWxzH5VrHSMjjpPOkK9xuZusCgq1CPFQkzE44
gRvD/Pf5rDqo+3+ebh/dC95ghehZaFO3LL4KuEsYdfjJD5YcSOMyMH8OpXQvM5TZtb4qVMc2qLSk
Rj3cmDb/GvMZc4o8lZW/UzUleue3utLZuL+hpMOY5hvu/YHqK2jxhtpmkpBr+8G9oAFfVHvSbjFU
zdwnd98OwOgdF2k5pdb13a1FKP0NVp98om1FE0QLBQu0WzUFWP0xRdYkeaJsE2Z8Hf+Rm+ViKGkN
8pSivu6b3GDQMiZgJj0YbKsFjr5jQEtLD/z3ABOT7aCDADTJKIxrRUIJh+8nVm+eH0r/jHNEvmax
MXyaGygbhV3Bj/aftZw8CWyFVFnHV7+dI6zRpX2wbObpjaJhBPSx3mSuUaNif+ED6FfHzEtO3stO
KCm6i6M91RKQ/za1lNUdnfwNiDowpe8l998EP8axGgigL/7XQc+7HQGakhOlFs7HOBz/V11KYBle
qkrb9g0dDFNhHhpm4nKPkb43vYXdDl9OpQiWzUD/uB32HXnOPXuwK2mjME0XMgt3GA1XONxrp9vs
NBBe0CfsOLuLD8+sFeZeqSmUpFl7wYvNg/iR9yalEbMWwEFnv0qU5ixMghty/NGiOSMfE1C2fr6M
HovQ0fHjQpOunSt/jBi9IHwcrUrtZZ3mlrYyIk63rsFbxcjsZn0uKsKoQ0D2/pE0u0EvfXwfW3LM
hy5TuFTtSxPdb1XesXG/WVPmj5aGnjOLV5I3wS/8Ux4yxr1aPVAR7eysvNOfh4L2E2iuNPCLyDEU
82r4TjCO2lxmGiKtFstqOFMmbvdfMmsApQWNiRtEoKx/b1+S05JSFu+iXB9dSQog6rcbPGb7fQ7I
waOoEoJBZNqzkyYdRvkbzcZfogJTUqFk4dzMh+EVsSSd+T8g263FKQa/DUcACzxQelH7yRRT2ryg
O8N/834C2qllaXvuWnMjBB3bQp0hqYrU4JDoM22dA6BtzPc4htSYp3mj8U9QtY5cfVdmZe7/O/V/
ubJXxs/h95gv1iOJSZyaUcKHs9TNd1jc4RMgMTAV5N3pTisDF/vXwDuLfSsh+ibQjJecAwy+WtG1
hawZ26NwTZB8S1IBd0PiZR8uCOK6Mox63SPXk3mZjDiDZQIfmSzcMNv6bd35ZX0e5ugtlwM7pVrh
y5pMgsRxjlvGl2PtOeAuXDNJ8hTX+KhVCrPl2T67s5aVgOrP/5Eip8kHjiTGcDXM50GP4w7+apJ8
2vEWv9Q/C5mTUnV/fo+JIxsKdG58O2qTe/zUlqiLsvT9tZEa23bh4EJxf3CGaWz9gRaPLZ0DD3px
5dk9JX5+up8s2d9OV1cITmUfOxBShJaE2KVHFAM/E0O0VlD38Zamlx/1OL2yVz3cH6rWIpqXQFi8
OoJSqhBkwkI/RGBsHUPn7mWD1M5f4pR8fMtOZYI0x9/cVPThGQ1mqhqm6aWMvXcjXGOKwJU+pouK
uj840pOKDJMMIVdzomuHfMNDLvozA5f6fg+DcPDxKDF4rgnsqovxCnZFG2wb5CWmu2kCelDlUk3n
GTr3cfZeXj+V4h5bJV5brmsoA2dtKttpEUWZy2UEFtGVUkz90+CMGU+lrs1OnGKLcSm1avnfRdtZ
rWGcRS6vu62vTTYxdxccYXOwJ8gKE5Uh8vJQydjqllaG8WB7sl6j97fZZ1XePbz+8uf5Y1TtncPf
WzQifcgOEx99nExVjdiWhPmz+gRNZVQx/nP3+1cbMH6wSCUXjGWEEDvMqTrKxXAZRTBK4SdgRVBC
fA29h2/5Tun+ne0ADrwvHYucGqxp5VRQFXsWzYKxahuZxmgv5X8QocXmrt+pu2H5dfBRAb0x+2jU
BDfbpTYkomSagO8NvtBMiVE4H/YxfxUwi7oypgUVwG2NlkWYlqMRAKbyqQdt9Gc3M1v/rbQCiemX
zHFxPYzqfgYWOxEqHhnlEOOyA5M1zO4wHyzM+V8PjcdMn9VGlLG8D/DGdg++waG3l4T5pICjHXFR
bCNjiT1PHk7fSnnY1PaE45D1xo5CVM7YUrhTqfYJH01DZSAFQk6t7Mib2Eh07lWHAuuNVRsTRYUL
uE8sP8d23rYiHTtZACla9FvXwmsDOEjg7luUwsZwpxreWJ8zjeE5SwnaQz+JVV0wHbw9zjYX7r4g
jyKgDMgPHaTDWxU1eoIVHlLaT2ATT0LtJSICA1s/v3qxXZQ5afXTzjpLJIVOFl5b1FBGwBpDFM+5
8iQfFVUhzq3kD4xnx+QA1M70Yf67NEGyBlAGYon3Kfv9TufYMtzvKbpliwg51YsCkqW/Jufmwtjk
OXAUn0B2jQWrwQ1LYun44Mw+EAFOLIsmQQGoLA2Kp9LXA4XN9vhSiFH4veGVqqc8mV0dqsANJXH/
J5AoYnv4r8DEG5f3ZCCt5coJI94AMcxrQaGpZ+BxRbYxq6453mZKkEgxRv7tksd+NfxM7PPEzfAS
/ScSj6Mp+kW5jghzeTXmLBwk4ig3rWWsdDHDoljIPhY8gyRUZ25WtjjwF0WHLJ+jsCBVPa+Athor
4th6vQB399GoGNe5844+T0U4rFFxQYV4doNtIw3PBDTemvqXIioC0drcEa20pkCL6C3Dky61BNIf
JLHuOyxopFlkjOiuihGbKLQRQEHeuY2v/P0imtxouiILUlWt24AFcDRmmM+mvc/JHEwmQmBxqCj+
A0gIQQCbDNg4llHHlOpVlel9X/ANUYk7VbHzuJifhb0GkMIM8NQAYuuYI0DO4sAJ6FXYThssTSTs
0DY3R010Y30WEnUGsYBY1J4wY+ONjV0LEz0IDhppbt0T9oHe+ERpsnAIxqZpVal/prWbt+SyhuRO
9ZmuNr58RPAufqURGwXKoS9zVp/2HFNv9ODJAZnlDaVurBaHWza6ChlOV6It7/J1q8OHv8RAvy44
tBjqlg6+RvXsWf6/Zw7BLsCbrJhckaIf+XXEDNtDoRTEEswyuqoSgBJ8M5mj+33BD3UB7P6mcXWz
AbJqTg5mxmznGdN10ryIysk/xqSU+kJDu8740UEifY6kIkrxby7s/L+t/yJzwpekqg1jq3oqUb2a
rt1X8hLBXANqNhza9E4LQkIDzH4kdl55m18AOLm3s+WfvZUUvQSjHszBEj421gu+3+NRZDhJmGaD
ndyNX8XimybTv+VlWGcjzxFoV8d1gUevigVzlGAJKbep+GkDH2rqt28TreFvEjnO1FV+v7BwOwEb
ILq9fw+2cXSNnaIgVV0O+BAyf/P2bbbC+d7xPFTZ8d1t/74/gvibM7JWNdE/NnGCeSfsahT2kVzE
71GEuNS2+EWM228WPA1iwr9Eec15XbtK+jSiet8adK9oXgLQZTdHgvCHMbykwV7z28ujeMwEJBen
alnsTByKZW3NhN1MbvJaRIgrY1HibdKIWGD74aiF6G1lsaorruc0DdPAydNTE2ECEe+zd2tZJVgK
eQ7w7QKD5OJsE/Tc6qPVuMa06A9JK3iNRz58clrgeJfPcFklv5bZMs7VCpnakVXrDp4woc2oqXHx
U+d9liuNY8TyC3etpBUAzxI599/wBUoJVgrv/O/fS/miIRr2YQU64pT14I5YCsuWk73v4ILKb7FT
PjZPLsiam8wc99duiD52YtsOtCd6dZq9hd1nTsWDRElG7MqehlkOv49xK/l+aZ9+nEdwSw+zDUsT
IRxYYMgIU/UAA9+T52FkUNjSXL01apogaPCA61qNK8THTWNhHuTrk0JOjJmBNOw5BT10l/nZvBT5
2BEiuboC/BZap7i7626FQzHPzRhHYy9DSWEbeiPKKG1hBgHe0uzoihnK+FjYBWlyt6U7RPE6WYcV
yEaWd88E1BZA2/bj6w/UT87bGYzSDnLLP3j3apnmaZDCmyBz8lZtLZvRIKQpKMpeP/8Avq99ASms
pbSWm7fg8TeFUpn801bSaPl+EsNNIhT/XnLwBILOs/USxhM81RGru0gEMYwJ5yfEF0R0vh2Ggnoz
2726EH8vKtBTEj00Mqmqo9qXq7fTM95Wy4njKaO4qcO5HnVWKO4UrMhDjH7jPPPS98T6Wwyrv2AO
XmEwcUz9jLfHqc2J1IiCknRkAjBRRBbYaeRtWQ5rshWiVCHr+u9xtyGtv8V7Gv8bIf2vgh9FWZ6u
7g44tiaXewEl61gaxcm4ZwGx5RQJliMkGr7eXlKQ4FMZ5cuimm8TkUNCYy7SR8m7evcpqP33kFSs
mTBdsAp4kvyoWthCAsfX4Yehzw14+8PaP44Jwoq3/t/fJUnnT4AOCVx+1Wri9TeLuuSvheNMKMlx
2UjPO0hB7ijK+S/T6xd9IWXPAjytRaf+0zzxHbWsvw5GGulQtwypmuVtRNOfGgcYd0SI9O6YxRD9
585r0iOCIwzOwCQt9YE0A9L6YUvDPqzm1Jo0HlDkKJDajXxun2dmJ+y5a6DPATL/zQCe42Szx2Xn
TpRZifpm2F/ZpevFm+hfokUaIVt72MeInfF0nUkjtX2yS/cWjryr2L494FVgMrYpmxnk2uKybeNY
FUx8TSoa8UPyE+dIVVIDsia26NKcoxNWIoxtV01tMONLFpPPrhcX7JNpVthP9vuSL8ywGoXn58QZ
OJfu+ueAN3jXidAn2mwfdxEn/yYRxF/uoCMynvKvJOxn/juj+20bMlp6sjr0rDRVAe5m5v6KNtJP
bjqvgkk8RsOvw7iSpL+IZu9uq45uHXRD4xs3mwvT03SnU4GRGYHHT0vnVrwqmtKmjuVquJaENi2h
muP6unE04nkib9wVqcr4xu93mpQFFLGVQk/7JbhxWJ/B9PBQSMUswhkJp9r4QVi1bLFMxdEZUgHR
STXjuijuBeq/eVFaOBNukZk/EeVHOa6RV8dBtotynDBDD2l2YrFDrFjsWijNdeny69JgWQl4++C/
wo45ujGhH8kRAjPymCDMoQ6NQBPqUNedoIxoS2ZwEgTPKs09b89cMVTxQoN293lB7+gjhod29qGS
geLuQJcDK5nh4URlYlro/KnmczfjALQu7YOhOyK3zS5+PzEJay92b2hdYY1pj0AuKRknv8b3TViY
M6/eOh7I+s8xuj0vMFGhKqmwC5TFlxLd8S2O28zwBhOCj0r0We2cMtLF0yKw6GXAZ2Qhr9higono
VggpMVX2H5b1aORqVaQtjryRE8NE+NR922/C5d3sSxzD5GZNO1ZtsrGgIFvPupbnHYSjTjJLlB+S
E1ieXy6+9dSD//GCgukeQJ3kfmaA9M7coEPmkzYJjahRDWd6SyyXVRLVfdzm2HqFZ86oPRAP7x7r
Dfx3OuqHv0QjD6+BL84+eDhi0jq3VkTTzB9VmpX5hnL3P4lKETzLMvN1Ka3dtmguK73IRnwO1wzn
Cj6M9bQCDKXjY+x58cx8yVOzHJQ+wei/ra5dDEC8/AOCuh4sBLvDR3cHB/vMZ6MD79V7VwBsPNuF
pPp3wbj5OnQAe7ByLlA8T/K5PUI9CMLZmRWNoEgicfi+PJ+w/iyyfKDa0OJIheYzCCstn4mAFv+0
RpQsvm+ecd2F3WpTJre4zHV4GnrhuO0sQYVYbgTypN74mr1CInpRVhuTw4re2Qyy38GYSpVaTqTq
h7FpmVLPVvzUT0QIlIwUv3uRnVcLab8cn6ITt1m7AIxViEChLgMbUIR6NaIs1j7HTfTZXRjIPiJG
cub1TVJS5meDZ0BoL6fgmJ3BlFpmP95z5+xpn2EaMj/XWr4/KcoXCDLk7gagcWrEtflJVeX58amS
XG8bcCrLypsTSBTV71AmU+q5BzoT3GqRbYvYrw91k55cQ/O5VW8Hw0CeUnmi3bAlFAyJ48VOg4Dt
iCXaouJdepnKxs/My3q+3NwbKztiNH7ly1DMaGIOuaCGiCt1XL+pdkNZ/cBpejkX+zC3+P+AY/Ne
p0MSHzAB2cFM6aN1j2TF0yHkMqnBSViy27TWUzIsnfYdNQr94yDRbEibRvMBQ4MkzAhmy+M83UOy
AZXO3MVGbEpvvE+lm6t4JyYqCBaL5FYL2gI9aJaQL674A4l0E4ht7NC/zlv7LMJvx9QjvpUs9s4l
qtb9gRNPtZGAnJOSX+a+o1Xsltv8oPEODaLxmv7mEB5jIhSi4rUaEnVBqHojs0VX59u2AVtLqRmV
DeWCnGtm7gTlWM1MNab3Ur6ydIcamtxdS3Fs6RkvZ/bHWdPQb1KvXtzTaK17vfTXLHjw25vF22t0
c2B6nCn9sltO+VrbliuWh4/FI3XvSFAmyLJBrWe5SuO40dACx/LSTwGTOfmRnh05sVaD0KrvqHWK
iJhurbPu/FdKKW44kEVtObES5mk1wwSOMUXcjp/m4zYCjnxhYnZD9a4OiQu1WAp0VBbItOGXrj66
+yqyjYtrPZRouG4nD7yH2NtpdI6MDer5C0pP6J6RUYNajZGDpBcb7U2OJG6bCgRQw5SW8Q50Je+J
2Ainz5sqEgQn/uw62IOyPDWRqIk1iTAFAaONsUQkxdcoSAbImStSuyow35c0l5x0p1z6DxCPTi60
qwzwuivh0tJGgBM4IZ68WAEwjwXUvGoiH2D1tHx/j4gjYjAjNpktv8gaICa48ta4wxHd2S8b2Ilp
kyfZyE2ffHu7J+kVIoW8tB1FmZjxNF6ZYUuTZZDNPeJ96iXt1zilOOHDLc6F9WEK9hsfspAeCP4o
4DkRLUKk1j8ASUhBkhBduoPThCJ6RbDaXt74gN8YblPWEwmyBibmYoYraZP3x8ZdlO1z2GeLe6/M
YB8dZt0TIxjJikU5fLKnrw35LIbp2gTBs0m6vMBueYyKOrFlDIpbYeTK3hRLDRFRQJvO/H8MOB16
R7yFD0BpakqUDmhZ/9OLbKqgFc1KiNsLjwB+We4osqDPeP5c3j+/D0OGL7kfS+k4bzIB7eMy2g5O
2hvLrNPo20C/lJW+UhBbZ7WajcFV7Qv/Im6cwv4i90HUVGO9wdGWytblqZlP4mAxM/rlJmjEwG9u
GOf8lY7LPktmDG7vdWjnaq7O/Pn6CJnxgBdDu+SWiW98Y/4MGYmYwGAzp8febeJvs7v9nq60CQQa
Grjb6c/WrxTkw6MQprYggxwp0sX+RtStIkKTqUA4FJ8vJGHKOBlaxqi8YbVgpq55MGJqaTzn1EXh
xWLrk4ZNVS69dl6mMTmRg9Hx05/zU2/lHLDt4dJA7dJmQpMKXbg1WfhGSS6Oyq6jPidBDrUEbGsY
3HTWe7vmOaS8h4+qzWD8IDZskuUO49c7lSmYY+5XMQ0at5H4IxVN0srBa9ZPNtdMHSsAndb8+d8Q
wOUN433c2IXp4u1rvjlYIcTsmADvCGUAHaIzIL5r0B6nXX2vlGCIEDNjWC+CH0cGXqQpeuknWHmS
hGK5WsA9kQx83Sm5dSN8RdsMsKxlNfcqVAvVH1UPM+sO3gBs3cYIcesh/Btp9gf51VFY02ATqUqL
4Qp51ZqU1ohq4MSMM58mqarwM5X8bVN1LcpTKl2t+oz2SUGKtj95PgXrFpYSDntFScap8k9FOQkZ
fX5kEiVe2wenkuEoWykBIfY+JqAbfqlxMAY4/mk1VE145BKfCwwP/6lLXZcSPgAJLB6gs9f9mW6g
wq29G95JxsK67sMXKEr5RuJ+DL3N2LEZ9q+Qta0DA+YOH7tt3d16u1DYgwx+hhr4tOkKnn5KZMBl
u+C5ygev7UW2pTDgq7RshO4ENOr4+6SGwFpeoM22PSU5C0GxNEd4HLWtg6VyhEOmUjRjvIyIRzwg
+aCp38HyiyEpjzOgllqxVCFIqjNQ8QsSvAV51CbfmgKpQmxl1AaeZoeIlvrEVdAPdlZqr26uOArI
ECRCNPQfAu1rRxDcvigQKNba4dDXsp3mEVLequ+mZi4j0UB9vfAyLoRunmlSe33+0lAUyisj7d4e
AtEwUZhzpagTT0nbFXLtYjxYzE63aujC4qPY0GBR27vYsf4xDFhesjeYhH6l9Ud+73nGl/ugVFMF
ZFBFnetz3U9qS/lf4nve8FEkEExCenPyCZItQodS+Cwmb9Tbq5YWEQ8Sp/raAaWwUOy3+WLYaPtA
IQdjn318hiK26/oNFFv8fxTDtkFu8PI473yBtETnLxYqViZDCT1N3LYKfU+1rlRk0DUsY4PJxDy4
f/lab+KkkACPxJyXtlLZO0xQCgQ4VgkK2xUV7JesACqL5549rATTjUyvYdn3gjbmq7IG+jPLK5/n
IDL38BsoNndhObBFE+OBjjoYJS+N29huKJ9xTBRIkancP5dvRqEvU05VnaqML5VErZT+pLiJnCBe
MFqCHGI98QEikth1rrOggfNwNiY2o5Ggn06a6fdLyZT9KrzNXvsJHZRPurQhUBililqgbITcLHyP
u666f67g2x0hFnDXRcee6+jFV3m4O/moxNW59im04IToWX4pndfeETLJd++EBOng5SuFW1aNY6Zm
SphFz7PiJ2jIk8UDvTzQ+89RZGc+I6hIrZ1yGcTdqC6CJ5zKlSe3En6jpRiV27jf9Tk7qhi3sz+T
8Oc3VPjbBIKJC1JzripdHbE588Q6HkuSn0j6i20BwY3pOriUpmuCp03qohkdHiXlQABY+4ny6IV6
1kHYOb7H/C5cVQnFt55rAhkApYIUcQujLKoWPXRzFq47wZn+CnLcfyZFLAQnBhvIq5IVuyFMeVbq
EK2YULvzHt+FgAEhRZK3xSV3AQZ2yIheWhLOfQOcrUDwlxuPv77dC6vSNlKMJoZnEbKZvWaO9RzB
x5ZNVWRJtKBnJLZ8iaLjicwcBSJ5jNQ9Wr9ykKXmhGAZeJMiDYzvqLi8wmOCk4Ne7+0ocLbwOFrz
F551HOGlmbsRCOygc2VyP1wYGNSyTdM5QOqoNUFBC8E7RsCPMzzwlfcC69n2qEdYjM3epnhemK8L
SLcDBHt51FBeyrVCAZev0KhT3ypKJ4OWMm1V+47AzQQiF6VMcIuztF25WLnlT3qkLki2HBapxQfI
yAnp2BQSdreXuCl+Knjjn4S7NE6gwp4a5twm2SoRI8s2uE3nYsZ6R7HVRAAip5zw/+IjDTDaTXe4
4aJ2IuZR5jY7+yFf35dkk0oZ5dK1T97p4ud8/7ftPATpSnmD/yp8cosxlnV5B6EuaEyUNSyfGyGZ
1p0yPJXbhy6vIEoqDltiryjCgsZbiAAO/GAQKJ4Ozb+v4MVBOOaZL25oQvNpDrfq28MjjrrP0kAU
k/ym4lAHWNcutjfEJZgevbSU5g8l0EZNhg4QKoIX3ck5X+kqWJWzff73nh0YjLdLQ+Aw18SBi/Mq
Thk/dBkfxcRmq0vUTTuD5/NaoxhUhY3PBswPAe8mGKFSu5e5Ssac0CAasBGF8eWr+vr3eR5KBTSq
oBgVCjiK8SUenUOfK7EC8jnIjZCakeBRw8PbXTsoo1u836mAyH/aPeu0rVCosP5q2QWRAYoNOMp9
HP2VQN3Z3HbhCfbXFG28dNIqyipxCtYWTKB0z6MToYFmMetdktxD3SeHmeVQDM4dhC2dOE7uB2Ye
Qsg/oXX7DaXwaH/UMAhdMH6ic5IjnsSLkEzhc4+Xof+yRRnVtEuqr9VwKOfJSBFQOR65CsB9HU4j
NKhG5VtPbictNsefp6XVKv4hACOjTRab6BYDS/3d9Rx4FE7Ul06YTJAlvmRkoy0kTeVJyQ/TfVEW
CZQqec80p7QP1YOK3ZeIxJTg69cVwJsYCjAyw39YpOp1QNeEVraHVp4rFDv8ghyfGGIgYaNVp3Rk
8bn8JC23+u34nBMWO8XCDEGf6RHfc8GUETKI8WS4FmvQ4YdjdOuBOtAEPnZjHt8pTWDB1DDfvFwE
vjpnhg9yU/aBV417e+Ube3e2hdnJHoTCoQ4dPeUT5v0ugEYHTFq+el75dlN+uuix0aN7U28IQE4+
kgiDy4OjRZNS3m4lZWXK6wYGmQNFDKtJEz+8/1TRLyBzTyfuMpl8OWpWDHyj+5xx4CesD0GB2Bye
L5aIRDtRTbVmNuzEJ42KIZ5TBmZxUruisUc0A7HpqrsxK+sjyVNklHX+doMsqaoPJ83+YN4LKbii
+Y8Z1BkQku4+AQIpCdZ0OK/HhM37VfTyBddd+sXy/dGzmqVYY3QsUyYA1+oiKX7s603srUeyrBcE
vEo/jGbt7aQYX72Ike1IkUE8oG8JbTb8lKm3G2y2py8e4TDSDEoRJI9GPkD26q1BO6sSnr9TI0Xx
zAfa7RL6hSdz/GoRpbLRWdtfBhDk24MHWYGKNkbwNdWv69WJFDb63yi1ZClT7xZJafh33T/koew+
FF7isTgP+pU7k7bSO5HvDk/pEaxN8Pnt1wTJJDGCTZMl/+EWSHFGZksN4YLURwtqNKeNHq7yRzif
r5+y94kBtddNceNNdL6YYk3V7nXrW5PNO2j2LIY00Eou82DJTvBkDed6USt3pef7lQ4mstPtpPtR
qjqed3JxjuWtTKVQvnR8iqfD09syX82KN4bhrYn6KHm7NIyx9htTxFAU9QELnrhiEZIpdGqRwvo9
S8bZA/h9F5c4rkD9IVvpIPr/lSilQvMDW9Q1XgPN+oq/oSwZoiWi6PfjylXZ6T0GDe7BlbjvS7ez
S0ap4Jp5pO1YXpSURJSIzgWfKYjxDjfpNvQmK2z5EmG9CpGNjYC9fkXfOO8OggLL4YUhFVDyJqb8
wR7nU84uaGSuhEGCdTlTbebKms+UOGuPAB27yVLInKZXMDcx7beay/Njo4/FXUYyUyus0mVVDWdz
NXEeGTckv4NDO0GvY0xM5VJ1j7Y2ivH+v8Sdk3TeKY2VcRdiOQjSQtf+azPdUjma4cqD5fnCRIsl
HBvqwbs0AiNT8f+YI0eNuUT4xJqaWZuBuJo2NBUueo6pHYAtBv7Dg5r34GSl89Vj2G4J8JSRKHzT
muGv6bMGYUSOY7DtLaAQ6/PNrVosXmUiDvxmLSHur55tIo0hv8pIrkm8g/klz8tDaNMqfD9oVLMP
b1U0qSL+dU+Hjz6Fe8u23ltuWilC/d2z7oZZq7DPJAlI5NXmKbdvPmKlKMbtoHUTNJC+lsRsiru+
1jDS1Fz5xBp+88wc7M5M+248pEIlVOIVMsYCk1NLoqM+eFxXmO0nGuc2MHiIY8MznXHAfGWbe1CB
Mf7qj2lLTSsLQ5VAQ+P1oDjwC5Q3rdwk43+sK3mqOWRJ+UypYxoscqDmqG3kVu/aY/YBiwwtTI6H
sjxBiwOejjeQt0XIClOhAEJNShCk1bwnjrfLUKcyYnx+lsrZZZhEVXBGXXFaDkISgF8crv9RviKW
UtFd9ehoEu+Rc6aOzhwWhjlvQYSWAs245Z7hOWOyWxf+JOrg5fibyH/a9b86zYwnpc2yaqfVlzRk
/2Kev2DQk8up9YMJQQyRGUslHTaWFb/g6e54wzZTVKeqS5X4ecfiO06hvQPaF/sC7klTpUjuLerc
EKHcqxchOa5r8E93Wj5PSHQJIJobJtMqxEAa+hW/8fk4IgdIOHHZfUOM2CSpr5J2vzT/W5h3LA4f
bTolDmM+ClNxo/2rg9LjOlamvmQQaa4FnTrWHCOh6SxR7h+3iiKzJD9RW6ZHtscZfpkztqZjYPLS
gRu+xAyFXtHsP+hyQvX5oX57LNCbAKqegkGksEoVm3Cq+7gGDSwMVABR1oKx8j335W8isoqv5EdI
Y5coB+7cvIx/AKJwMR7bKb2lTsXtJ0crwdMHRTEhjj5Iu9c3OMskWTo2zHHNQv6MhO/24PiuOFvK
68OLk0YAlm3rCc7k4HczHhUDqIftmSelreliudwi19zJ6UbW+ZJ3Y9CqYigzkVECRW7x+8xd0So4
MSI5STpbKq2VzUfJ7X5AkNWvY39Pe1SKet+qUZ0/PnPb2Zg6gnk/KBYQQASjPsJa+XGMcRD4CNcA
CItH3jDWgkuVIl0ZySDT9yU+BNyNMJRDjdmk/Re7C0K97RBQ1mCt3tV/t1GSYwzo9pP5fe4c+L0v
Vjw7B6lapsHJnBk3SlMSqavS8Yzawp1/g7N8ilmGTGRA/z1RxBvRKy5+DmW/nJiDvHFx/6NbWidp
Nd2kw0ONulnaUiZ3ZWyavQMMN5rHxifjlUIzlXw9+3ZMSeGn0JzLdvFmNEdG2/xTzsr+FKIxNGNU
hoIlDwd/OMqMxBHA4fU0cbvz2tSY1TR7f1JkTlns+1/SqfUTVDJyKZPCg75Vaqvp9sVNLj2v7X6D
FoLP6xDQ3Yv7pSXiee01CQkEVV/elN9Uz2Q0vHKlFjg0cJXdJxOxb0xeObop+LLVX3qNSPWYcRsf
RHSlyXDOhU0fH2o4Px5smRS2DxKOlIOePijVdq9NwhO+vAMBva27fV+BLfPtyishSiY89vRwpMtx
X/ylVy36boOCSX098cqnr45mb4QjCrbZE8jXBuVzvmIuW8/yz1VD2ywAPawmML0PkKd4Mpks46tp
Z12012QKspIujhA9RIv3xUkVYgNy4cGGBJo83yvsrDLgzl2Y4/174FDBFQzpsju+j7tS1+S5a/ZW
ki2YTqmuvcnlXc0c/ErZX6AZ86fTnqyqN6f7abYiCfNp9LMPkCSJML9sGQnNCk1+xWTx+7JU5UNz
GREgCbbWs7GC91CNRMfMvrIAYo6hBE65bIH4tmmT5ntNfC5yei3Ugw++R3fhe/bH+4rqhSxUqs/x
II7MpNpfs/FREtT0wQhxCHmkP6vLqkRLZ8Fj4uOvX0JAE3buY94KQrMKaDVFO03YrqX/UaWh9iNy
3VpSvhj0w1JwWnVdwCirKUlQJYjllgxpx/szVfUO0cA2hIqTV0bDqqsYm08gFwjMupbORssuU8bO
LoBGwfQqNTUIpU8Orw7h3FYpNnB4aOHe+8Iw9cMlD2Ko+Hnb/q5CDlzdovINljBBP/HSdUTi3xtT
1OgiZR8m05ccD+WNVok4eZznSHISUMjrU0hDkyqvH/v52zPepPxgqho7ERKykIrwRUp/oeLhaIUC
6N/ZyVPJR4k3EL5dSn+sq2mgLjKgCUa1IhLg+Qm8PfJg8l0aB9CLgPMNtR04NOReyUHQgKwuA6FP
r6+oRqaFNUvRP139GqNq1iSHnV2rx+cuS2W24Ari9BKEc+iPGi8qT1pF6mM1C49cT1WzHaj+1QE4
5AB+z+vZVuq/S3G32SSDqeKLE1cR9uCU/xSKUORoJikz7y4mdmo/2HHROYOFxcGZFlhiqz1zyaIj
ofaINlIuMgYGvNzS5rxqcF7htovf9q73ri+zaqRooc37zDBUyG+VpLi2fn+c/5uV4XX8sFWjIenY
Nd+zcCUVwxZFLcW3i2jjtEtrcNj/whALEDPrc1/RDtE7SqL0FIEIxomNQJvrI6wSg6VnJOGS+eJ3
DQ0dfh1Mf6mRrQevragxPnszxqvxL2soBf8Umk0PHt3boNQ5Ytj1UjfZiJ3KsLRmtAQUr8nCJhkQ
fYEHGckcuAy58PV+lKGqFpkjc6cRcV+wUGb8+SmBTCqbSg52hMPtsssJghmm1Ry81+bS4SInzwFl
iBLIuLX+F9XuBrJUcyq/XBQ9/MWGP77WkEfFLxw1SmqftqnzuEZnMre0wCiKYqkW8agdnCKgI7R/
dZ9DnVvWivl6QpcdxRPzb2F54J8Msw2nV8NKhU8RyD9UTE7UxHVOAc91v24BL42GSqf0vZzHRy8K
cHqpQjjwraGfAafIPIbAAkCGMzYkMHmAWH9VVWdjC1vTFvxVMJi7rsRYsT9Ogd8z3WjR5MQgcK7q
UKguHeSR/I3PgdjKRpM9EyaCsvrgZkCEl+MwVcXR1BVkMPysujpnLTlpAvgxfMZZtwLw1EGcvHP/
wYOxV4OC3LzFpV5UUvksOWUKaBBro4jV3t27zNCN2QagN9frQoXmiO7fdszg6hH6He4TQZx1rZmg
8iZeWLFFhXft+a92osN+SyK/jaloXXJPuvmI0sLn7qgeQMMZ1HhTRrq8RPub0ULx1PcKcnzEfE+7
NsWNWge6o27oCO+Yf6yzGxq561/dNTRlG4XNzkHEu11o3/HCcz+uV8cinPDQ9YeL6kYvzUIuGUcX
Ik0yrRJgxByCM+De8Yq6FsU4tVVpJFjYZSbLI7tfAuZzvijhZeXSCWSLl4sRfORJM3CNGKeOrW3+
kzZockgVPY6vv1TlvWV+COvzuEXXfzLnEa02WUTrMTSaygA8PZszSyIn4jxBdzDn6HZ3SipQIavA
FrsG+hVNZdjqCIOgzKDid5NtigFiwBSDKUcq5Z5GjMT87Z/Ht3L1LmX+k8WfUxBxXeT+i3ipObzB
4JIveCH0haIDw8AWUyUsLB2nutZGg8/a0dtJH2oz7mVcEpXnaCNLpjZ79LhwL07mWiQSeW+BcSxw
9hcPmeYMpsSAhsieD6tNygV2lHrjhdE8d60wLguQuCLywTSNsKZ8Zcsmgc1fL5ZJ8y4u9NnG1KcD
UYeprMH7LU1k25zRJcv5Se+qt2vnqXEgPK67fv4BMhx5+c4Ab5THh49xbcRC+lKY1e0g9QO7j3qs
NNXoJsdjZlDrMtmzPwev1jxuJQkZc7mgJcU4XiX4UCfISEEB8pJRSBSZnIlZbnhbdAjuUIXpwq5+
amPojPjG0S+FhtindbSiRq+z6KuH7huvdzzk4/uSNUCAmDDoKuGRk+dOBHfJcPC842FQafxCFMGu
2LEvFrPkiSKrpqChlUMJDTDTnv6hp1kBm5HfWPpX36wKy8Jxe5wGGiAcwA4UnMKj+ZUS1UQAo2Nt
lgg1ect0bMd25YTFbdEjaGOZ/pjweR1VxZL6O3kf07OAyEJD3hYjT8GAyO3bQohgDJDIKKWXOFGD
GnOLwwQnV3ewYdNslDhyb9qaUtCKdzQ8Ktrynj+mL4cEMzXBucGQcM57BUs/LBs3jLJ9WCHJpMT6
5MmY+meQTPbEhfLjap0m1gYbaC8Q0rZQqqS+bocPU6tE+tPfhn7QHCLOmuw/1dKTbjFZzPlh82cD
PWuAat0ZDFv96AO0t4+914/lJt8Gr0fWuhyes210mVkANH8NWVWHEpy8TW5lZC7DQa6jN2ycqlDT
cov/lEJex/0N6vXeflMSane4+sjFvbDXF0M9QZzFoV7ONvYprBY3EVWuKHXLdjTUsnJziGznb3o2
CCiOZEGijzg+kZiiy/c3sso5nVtoXq4KOijl+K2yjFOgCIs/DWlip5VB+LuJtoiw6vcMlc29u9Z/
wGBobAMr+mE+Po9QZzJliRfvn9/7qkDnowwk2tlbRNfJAex/w98b5GvkZLJ36aSn4uwLcdLWiqot
2ud4w4oSfx9iB90nGJ4SEsA+PEL66TAqbMk7SIy1pgbd/bVHsXPri7OomtFcpfj6WN3VJzBCob6n
B1e2kfG/OCuzGCvNjLQo5uBIg4w30a1wmT0vtezD4AqXr53mLJBHSeMRd2eThrMmL9Q/Zhp8NDC+
bA+q2vCI/sqYf/DXhA7zOPBUWFZN2FiuS7huMqFQ5o8GUoqWjit0DICq0QVc+fJEOn6CnDZ62igl
MtyfSQMreizphsP4gSMgz6/XHA9dpn/kZOOHVp09s/GaNO6gRQ0FlY9BkF/jWhKtfqsAZzok+VT7
ELtTM5KzW5TkgKN9MS4rKXHZCR05zS63PljQnjp+TqexZZlPB4xackMGUH6qBTHkXiRzb6mLI1Va
7CUKOtofZ8yaFCqzjbOA0G0OzTb5qymF/CiqBgF51RY+g7ML5oMN1cLxZ9DxgihTFAJp0lvG3vUF
QIr8IlE/8ratm39Lxp++9PiBOLKrrk7BhEZnhou0i/gi0drDkdPTgKBQxlaGKeiEiBpg87zekPKb
qv3V6KAR+ICY9yCdK5h3mlf+1+VI54YQ5JR+TJH689T4WP6z6uOo3Yd8Nm68hF053lRgolEUe1Lc
9c/Mw85A99+9c8mnsfWHMu8nrFHmIcaIho3CgRd2nsYnZpswz5rs9lECJ3rZoZwTYKdabBBoWy06
rvXdSianh5N3a/ukszDZzl5vDn/VnJorUOKTaVoEP/ctVBk2bi1Gp6zcydKbV4WdMiiDC9kC+K1Q
IqUvazXuyvfmYyveB6wg2f6wqUdvR9AYlSttFwN25AARagH8yzWyuFiOVyg1jimUy29YaWnCAdoe
txtw3X4PZTEDwNZav6dzWEDVUrkt0GW5TXwadAPXV3VwaOYQvUdrVdSUxngS365vYYxp4tgfudBy
Tjuxoxrfk9WtoEzEszhHFgn/X/yHLZsQE3urIZJu/eYYxFC303e6OHrGIophKURMyOkkRyXjnamR
UlECXPQv1diJgzWDQC/y8kujoS1Q31VPqLp9BO8jK89pgBTSXTZHgXmQ8xzV1IVo8QRHOUsPkYGk
wrHPUKyfUl++UATdRhZ7nDnBTqrgbNiUcqebQK9XyNEJys6fYgw9jHdFoL/WWmh4GdhQtvIZtJ2V
ivikdqDYBuLuMc/FjnP7LNXeHDynuX1EKEmKa4xJKXSdrMO/wyiRCESqmqvgurmhmMupWXM2iccj
+kqchKC5sra4kKQCtAS/am0t+0WjBelpkWcXASuXcpyhjyaasG8SJkZnG/OF+SirzkTXaH8N+4BC
DSCrNGMesbl5Y64wS2KX1aCetdkM5Kyn8+9Clhkem2pqJzHx3byiBIx3y3yLwr97cxTxJCM+WHzS
RJzuzYVVIk9gi0Rl+aPWz3N08DE10WItu/YMVdBG49vsIDNi58qf7wNVzrQ60uQ8bUpcwJ27vHw1
B3KkwL976Lge2TiGaNKsgflr7UYnxIrXBQ7VGWEOR5eSVMuSAKJTarjMmTqlPZr9HgkUnIKnY8DD
c1DtfdhJVodL6UttjfgjODKlygrrFsLHhgxPv5czMazFsgPFmKnSrinQcmdhVt9k45xDHXQpaC4Z
i9+/sGowuR+N19mbcQ0vTf7LFbug9KnYnZlVbOClVcCfeyadtEhBjMCEpB4lJYG0XA2DqiGPuTwE
XyHQDyJ1S3B/7iGxeZRrkpTZQKrewlO2kqJXWDiYVa9FRobnhGXYBYyeByLLcRiYyt73oNyfWUfL
dXlfJCwUKq4Be60S/+jbBZwIHInkYGYwcFn5I5phGKo6I3p94RoNBWwYyAl8ap95cOUYb9scb9Hh
V5zDKKHokzFrMMuBstioYCWBX1Yi/4Iq7SVALBNwoaExBMS8onQBUtxEwjLB98V/s5K1C7Tj4fCR
s9xfVC7qPcuNsS7cPDx8RB6Hpv7UMMd80mzbn1iCs62+bAT9JgWCHGeTO4LL6DdAnVHZlPvcRUIp
mAjB+b6UFx2fAf631RnDlhxOAJCHO81l2bvdu4a5OU9XR5HT5OInVYlnP7fW9ohDdQ1bY4X0V1+9
Vy5hYNdXtl91AKOJ1qGCyIMoCrC38pVOBlfE0WiXCjcUSEF6uFpv3fx64wq92ih2CAlcXJeP167m
sC4G1kpfIRVi6lDPG1DTX3vUEiDRsLAOHZKUnhsZWU/QtNKoKXxo9S+M8wwCqOFhGqana/sjI3CO
fFFtYH4tyRq74wAzNwu4Fbujr0wZSqtAsNFl3Sboyv393CDfQR1DkIOalWigIxMV9SlAa4n/wg6u
C3UFh+SG+7K4HTYka2gWMagBDmdlnqLV1vkhcx+mGc0/3I+HurZdkBKkeprHuk76IHGoLCPHCmSQ
gDkyIcc5qBUhPlk8vSgQiIhr6TuIK3BwwudlW8VPS80lyjD6t1zBlFepU/vsmc4o/jKPAlNEZvmu
04fUnfAErM3z8GgE0477hOV2oun8Q9DhgkeAGW0aj/+i9kLLTSR3SBZnNXPlfl2X6JJTnJXTDtX4
LtgPjWDCDjLUIfqXb/MDDH23Y9GEhBYFFZ1gfYSdp6frQvy/hGH/jPHi983XKkrKaOTFtiuLWC7K
LVvgtEDjZiAuRcazt8xOodbEGK5RzowzI/tezABAUAnz5Ns6GMFcJsZ2C58a9rc4DooGh9oNB0Mm
69g1iYe1uJp02TnqPicsHQbbXaXJHcH+xCoqU/lzbHLI96iJqq+i5HlKCJxu/T51qDS/EGV7HXQD
EgHkJVkRKoNeC6T3owJZre2JuZ7sMYKurwpBCz1SkpDan2d1zfJ9AsJkwpYsFgvO7v75uTLP0ZOe
mdVt5LZzOM+I1g5/It+KkR+FAwxekUzrRh57kbL+St8d88/A6ACzm8g6bbZzS54ZpNzGxgMNSoFB
D2D9/TyTzvCGFuADeeil+wkVnS0X2FXXKRlmkvfJIA45TpfSv8/2RzbgxxMFjcIBk5kEccLQyxTo
7Y6NCro32GHWQmIbvgd7lDx0SOlV1ALS6jtMT7iBzbgzfhSCOMvwZUKK9MhUxotZ7rHC3mCCSd3m
n0l4R+Yr/btxbShyOK6Zlyx/ZFDWNI2T0XbM6r4L13BL6AXkjCd4W7ZpXHYMCn6HN1N8DhD5AcSS
bZriilJRnnvdZ12aC0hvIKD50sqyR+LC31KpZRucXdlm4KVcRw1fai+r/hzKRQG30jqzemUac2A5
PY2aMr9qygpnMCmHnhGKGzOFeMDNLzkFgSkk1mrrXcvl4mXCJN7moZGvaXtBcskatF8xmJs6Xfml
gfv8t1KchNADHBsKcLpbeVB2jfQaK/Npa7vkkvQg6rR34Mm0Q3k6riQBmFz9lUhbVbkQI55OFHs5
WsL3zInvyhtEDlB+vwsyisiikhI7VHWIcCZB1B8X09DStHDNakXOlXKoYGUfj8Fau2ywMrnX3+3L
LOxiPNWho86H9xN7m7tBMNoA1R6B/MSEbxNbGVrpuSNv1UxKQdhstMXUEYOIMLHrghyPHxefcXzw
LyyfBr5jZ/NCjusiWtw2Kv31032KzjRkSaRMXE2RJYby2juKrVcRv7KoW3c1AMoegNClcm7AKJXi
Yj17flLLV7ysR3WNcpgdVkOsov78a+SFk58wDSerm8z69EpmdqOfYT7wsbwfSKzC7OZJOzeZmqRX
liBwNCD37FMiftMhZt9rv6uLFsKTLvITrFbRKW+F+wghrnUYKAdzPQgH1JL25C2BPE7tf+z6i+oA
XYsohWh/LBOpqv8Za/vZOwN6eJaoRGl9e1M5IJhxtRDtPWBOQ9Bz5Dnsqfa7XrwZ641QKTJFYjjM
6+WZjyeKNnUVOmjawDw+l3TWzYoJpsN4pZyJgslYJR6T/QetL+TNE1eIYkjCpQ3P8QCQI7DCcCnr
4fJP6gbSIB26qym4u/5XbWSFfYIh34H+pJLGBkS5wlrJgLOXAIA3s319wHbp/hR7Q3F+IomRpsAZ
6a7fnrs48C27XPW0/sZoygHvuLmCpJAmEA62ijyQwHzw2NKdLtfu+hm6gqYFWWhhpWe1wUBVUZt+
xXqnV/rNcDh9nW/7U4vTiY3hmKV+C5snhDFqnS5MnF2LUf+eB9wLusDmuq0kejTSaYw1T58nE05P
q2lGrZWhxV/xZL1BdcqcbAn/AXMAO85rSGkf/Ab2fG5G3vLLxaFhqoe7Q4VR67xLmnW3nJObEoNh
wDmQKYeXrE3OSHuEmm2KyPcb0CrM6D0gdSDgLB/TEmC5DMXZH9VYYuuPTtkhHDWMHLQxF1Y/thWU
sota4W7ifogajvP4XvCTqxmeoE4cMwDX1D0PryoDteG232WrnuVYe6OWaZD6N8xp7vJYIlWSUTHv
eiuCU45w0mTs/Y2xTzZWLv06NAlxEHNpUuXFsqtW11Gn0DxocYs553q8gkjou24THsIuYpY4DUHc
QBRrdFJ7S1d8GzVxACSy45Ep/Nf3un4eeEygOz9dXg65gV+aXI4LeXdcUIggq18u3omEr6yfQz67
H1TDTetMAUFAMiVm4/9nb0VXiVd1eqO1lQJy+tD4WHp8nbe4F4RfAg64xBcN/SgnTeOkfR/HFCb7
ijRnm36e4CzBJeFrhxNeyTTqu8uettrAD+ENdZfkVFCxohqfjP+biak1I/1mHG5mosUjepaYLyZ/
IJ3VhX+rdZArmFzBkKL6UU+Qayv6wcNj6JA5Hd1ZSmfa4pi9JdVWHrhOtsdUJYOLq+CBLL5YH0vv
R/WXAtLdP5kbyiFf0VcweLjudD191+gE9dsuAyhn89ZdbaS7oJ158l2OPaQtaVcV1XINM1zzgJ5w
ooeDpCz1F7b+9I7jJ4H/g3zGITdKIzXRWCw/K6nNQw/kfb5cuNIbFBy/csZLHsT0kNDELrfr4m3i
4HmzfIcSscW76nm9gm7grir3qszU8H2ZUP191CGzqngdNAJvi+OvisIIcfo4HwC5h/Zsnw/s3sTy
q/hIVD9CrvyWf6qyRo21ZJ4V63ERow88t4hJRGCyZpptaPeaNR/NiF/Jrw9NdbsRUcrX3Cn/TW7b
iutDoK8dNjAGO1pesIeOT94cNrGxJAUghGnk3L4+ky0dkIkHUshHgbHNaqQR6NNEoobsrS+RN8YO
zJIsLwF1pgYoY9S+hySXkoZKV73roHP9uHAmf8Fry0rl91CmtdSVSyvNhSXuxvh4dMbr2/wGpkIU
0kcpDuMYHVSnaGvxDkWn0S3xU3QeT9F4eM7W/eCQtxdBycJvTXaz7OBGwrizzUlumsblmq7R8iQS
XMMqiHr4YgTXuKdGuMO5aDvEQ37VQpYjphdUe9kDPoxaoqEo3lhhqLdqqaiLVT9OutcLHsE7TQRg
ORcfNA/CwJZTmyxFttiYImIkgbNnDb2prEaGj+qbG0ii7t0WgSgtuJ1BGMx/ORvIXPAaW4BsoSpK
UDR50XUzYsUIqGkxiE3NOaVqvHA/fv49U8l6q2USfHZCnrN/76oeJqJcXkHskmq15EBthL+M5hA+
UZBYqMV05TYs4vjJrawjT5X+ywsmR90ZxU4xL2a3M+TzwbRjWCMzsWNUQnBmNrCJ4AVJDZKIncuk
MhxF7mvDrbNFMwiPMGSRVANKhZBQceiUgXQXKT7krK6I/3U1wgcDXlNsb9VJsvMJtl8aKIhbpi+O
vAf6/U7AGVorC2iGCJYo373Vr3XhxXQJkhqjagm/jUm12yIE5AYtiL4XMxKnusTeH10cKD07Rg5t
pIN2LSS9a+cbET30PVQjmlB3gmi4I0YEM9r3t5LqYhsatZer+qIxli2PRofMHLYkzFQzQ2ewJb+Q
xLLau8xQ9P7Aikp4VdkY4QHT7ErTQ5RUQ8ShzfD9a7KBJl/AB1OVyG+DlLZIoWI9Cv8BSwVxBVsv
r+IFCmynGGvYl5OEB1BU0D1bapq/wSjwuZU7U7xLAGMv7NHv2p0a56XfQ/Fd6JPuF/nYi9i5gVwp
qun/D5Rvl7onHD7yVxDjGZ7FsLezce2iO55oYo2QztLGQ+fLFzJyzUakGCzeOJ0SuvWbX5c/xQnB
3XidUxzWnUqVK+DjdDxlEPF6LX/M8JkZAs65gOyymfd4jojbfaEqkQhzub1ihp3kyQ2Hrgd8OUWJ
7Q/7uFOtc0kTtNZKZrVgb7qEkyve2za58ydTEQNtu6efhEcfM1pTxlfyZ9e16+vMppTejGz/fU4/
4//aJkXvp+mXRTIhfU+WmFjiOfjwOKo5Dc+PZ7gePJPDYdnuwerifSY+HS+YPSxuvCcDtyXDLlv1
GhRNa67aorAGgdqfQtlJfw8AS7ELZFoKDtJkurEZ9I6igA/FbLKfJIry2ePQf3Nnv2ljgNirm2vy
F/I1uGW8qFaCXDygNebLJbneUPn81A0FMaAgGnh73KBq4hEDE4yYTeVMsxaMJeS52G36C9E9z0nP
MhwPfPX10wPutEzlFHhg893DQFLd4bt4ltW6Lqk/4IqMwMa7zj7785VE9gqE6DUjWZMDEFAWlUGx
0wA9E1lPsw8MTZRec6p56xEaji+HAtiHyXXS6jXKr0QdloRNHZp1ysuUM0rdD1Tzbi569a8ro2Jg
pe/RhDNubFhiX91m4htqp504MLDysFWgRpJ87t4d9RmtaMNufinqAqKqEwBbfn6oEea4tKXw485G
OYTq6lS107axc/1nxxzwyRf3pr5vKTLlRKPj+fsG+iTC8jb2WT9dKkMk+lZnncaqOLcFguKM/V/8
VR8hUp2LnHC/VAMJKbibzl1GDpE0asgLr6/45R5R0uJYYO1eKyJ7r419/uiCs6TgR2nf5/fp4AP0
otAnVrGHcctc02yra5CkLOAfpb0ZZt4BIbPhaddXUyQ323zOlkRHIdZTQgPQBTPQek4hhxCnwZyv
TwSm8YQZzgC9RIOxq1gBD/IBI+SMmrB5EBsOAg2IEEKrXr5/33pS+xlmysJyL9HrOI1875/+V1/u
e95KtZtwyTujpginT1gOk5wU4L+JTvytQmHimHVXwClEReUMYbF6r9Aczn3gZolC+5PSr3NooJqc
dqqI0/AdhdYl2Mma6O2BUY1zxETQ7HivDiGEzCj5bVOMFg5IlJ/il91di1EFbv98oj5HYt2ZI0hD
fHIdhxgEDAlCe2HhZFtk+ynwptYl/OmMw67aNJm9R4Ff78eJXH9MCSqXDCndaDMXyqyPhsJ1nXAp
za09Ks2kPLjYXncCxKlsvxHJfmuGPJG6QBeLUdcgdBIIA9f+qC2tUmK/u3/jm5nABvfJqVYSJ8q0
ELHu4V0hKcRlJ2BzVQvGFeCCCox03FyWvVzveMNEuuJB3mZpYi/xEviXQySAHNMvjaThkoivpwk9
ORoUxH0/yio/CL7s+uHswUPr4PASE1oZ7yZTZuMEv6gnzgl2T/69V6x//jOlIlx/NRglIGn9BsPb
u8wCvgFZlFzvUC7eEDH8TsRzbI4mUUn/hjEWL46FYGQ3xQybBhbjIxk+hM6XAx1dTG54opZhG1Mx
GRuEt23AGriqjKImtJK4rF4Rt18IZXzjmi6r6s3cvOm6duyZHcNgPlWTiA0ZYi72TjoZechvGLZO
AzJrQY72YrRpL1HrpBaPUefbEpSfaXGiKZ1juq73in212RG3hpIJNokikvf7ozdWXUBN1dsg0pr0
QNE2bJedfIyC+vsSqXMLl6LIOmMY3iakZciz5wc54HfuO8EHVmMk7zrNhFbclyfwG+Ib5bLTJOHk
thVeCq9msanRSm+cOT5V7IgTCDXLYRlqy/P/nBNijYQFoSolWtuMcCipASYRzjUQC/ivK/f9UP0P
iszKVMpyDsY5pPX0ZvrZkbc1XC+IK06vZRXF/tYabSg6pr2hVz8F4Wsnu2lS0AlN+gylRwh0rKHD
ooj6S1mp67DYKNU01rrUhCb4z4k0J99PmQqi7QDnxBcLKEA5JP4xMM3qkDnd/uMO99Rd68ePyEQm
H/TFne7mpONKtUxSGvo7Yc+krdRhhlJO52U0oeAyr4slc1KIeXTAUSEKSnbrG0UUwhjSApyazhU3
8qKspElGNwc0MElqIio4cxJBdL2zPEVSeddmI8gS2ee90S345ndODORl9Kpzll4jAMNBTZigp48b
8BtpQb9+E+j2/jv5nHDUK5Ik+qp/V9pEClj+Bdqak1S4T+S1nL8OsK8GEvihZVdhNDLKOUDKjetw
icdo3bGA28dzQMB7Y6y9/aDJvVhm0Wq4CS2SnxvdnWCfpLj0V8dr+r6Eb8wN6+FgWCR2cCS4UL2s
AxlZYk5QmzXHvxi+oeh/ID+/695BcNw3VFYNjYc6M4UZj9pI+EEDbad7SXJMEYf9atQTrrsCJkil
SeAOedyg3e9HJDvq00D3/ae+5ybsBKnpMoh8cq6ItgpzxOyVByFQEVbOvZ/j0Bzvs4nbTx5OndP4
1EWZrtA5xwZvEF40T+eWcIxx7DY4NvYKeTxWrbZC72meDS4CiwDwAg3WWIncOYEAcy+PQMoqG30u
98DkfgbL4p4spd+qcpaPquz4EOSgpmuIEzxMxOt5XwAuB2kiOE8jOt/RxArpcgpLXn4YzLThd3dP
xqhWA2JIn8zsBR9cNO/zdQu0sqYhWZYQRhZFb9T56tgYOga4BS4wWFtwhILg6BLP2RRY/3aGA9/w
uVyP2j9q+PjzAfu0Tpu8yQ/ZiO7OCAlHXUq1rMUATwMRVGFUM4/85OG9xijPxqbm0Hv9Lv8gdinM
d3fFor+isIyXRpVCBXxzBUKcbh00accEi18WM4/Exq5kepSYKl7Bi6s9WHJTldFaYskemQpqnyDp
lujDNWyIphILqboZ4x/ZHAp6FTWeJPfrTOIlRMC2XrZiP8JaN8259O+iYx1T52f2aQRqSmUPgqlF
s/PJWnvnxfGm5Qr0UmrDEqwrsrTbERuk2pup5939ZEzmR7WX9DMug+3Lk+y0yG1D/90twn9C94pv
D7dK1RdFDHwDAjUWlxXCVm5zpO0cwUX+NlGzkESeA9sLT2eFN9+vt6Tyi66FrgFmE5dOvDpvgElV
hgY+lL5BmsoT5b7FaEf7bHeTW+zyYld6RzjIPPKx4/8cvK3Av657KFmRn/3yrP+AHptp3uhsqVUn
3kKzJLAAiIcYMA0qIqmf46LwJmTM1+5RtcVpHy8P2pePL9K7srLDqjjq+K7tCcfijVukDFLFXIn+
wjWCF7z2yAqhC2uazYTPOVvgJMM6KOaIwgtEUizHjjP7+mEJUyLIw6FFEM0cDUIjFplh04PC+m/n
ABVtJ+cEnOjscKld3vH3W8OL77Cf6kKCVJJGiaPs857ptUw31BUL2ZvRFWH6EaF9huc+G13zVi7p
y8fVikrl/rm8sDyFkRGJyXfNYrZdnWUU1ZXVt4dXBEZu7udLTfnqPZy1wT0P0l2dbsoi9yHPvM1m
GiU0ZH3AdEA1tW0q2/AdJaMoeQaznS/PfYQva+oW/Cm6n0Z6SvvMT4TTdeFA++rAuDUv9q1wYpl+
EvQNkEZvDhslaEv3DA2278D4REcFKJIkKZlBMzcLfUfkJxNWMpu6lWU+HqZM4TAgocIkdV1E1ews
UxavdMNFUctyDMZkVx4cddBrrwlNLmdn1Kih5FHt1i93gqTpd8fTCg5fwv3AsDtM45SL0dpG/4ib
C9Ca3rBORbU76wCq20J6V4gd/iNvwMQLYaXWk2n/zF1Jw3Kqkea/Yxx5XlL1HexD37a0s7u3aeei
2GXap5IrrG74FsdjU4uulKWsJIFDGxNG+u6Iiw8r4VVBn0zUcgwYqG48rdFZvVhQKkzQ4vAdcN0X
4Z7VR7AnDv/5lFVixSw1pvuSHasI0450LoRKzLyUYoSc/LDWkHHacvM7IgPMc/JRiex5cYCeO5wg
8zQryL/Fi5FEiVkypTMgOyELjUqPHBw3kR6RGCMImEVCeDqcJA7PHoiF3/pQzpM6u6YrPZ6xD+MQ
4/grS0Sbr8C1a9i4gHMT9CJ1mTh6ZY4qQzqdknKzo06ZuMzb5sQNZSFJo+ls08OsddK2+4XuHxaF
wI4BwgVmSUnLKA38DOu3mcST0Gojxgw8watcezpy/aWQYvC2jDCbqB2iNPiMjJv4YZuN1BSmixT7
MiMy/JNFUfVGr7JQT+ntT5AaCI8CPSR+9VwgdNzJwP2HlCtlOSuZxWH/9zEE3YEojRNcOMk4gxHY
3/ajrXHT8F9qX7tlEgd/lfEYmqgZ+PmsPStlVF8VAfCF7BSuzm5LpIqjkKz2UdLjYYMxEN/Tyydl
Wxe2OOOnGDnQ1xwjyXap53MRnp0LyitzJJ4Efh1m/jLHfwEi1g3z4r85DLqv0C6v2G6KOmJk0U0z
kZpr6zsZhZFQ9oRoiAZZ1vsFlheGBMqmNpGvPwhRLXkwCbXuZtqpDKZ7z+G0GZr0+LZrT5+MYgtj
/XkbWd50zeXMpgOD5lA3oAaas93qlzrXoysMBGAkuTdvWR+3dbDGPrdhfXminV18IrVEC/sdTtEr
7MsKdkF9p/P0kXzuI+Vyo/NDOIEzj55jYLtNkubdcOuKRToZTllilAQl9tD9qtWklZ1uJ+BnSpBK
aB+nMCzGXvRI6NCPQBd35jMwYmddX96L5rQkzdhU5u7LazrFE9ogMsIkQXEltFksTsBjnccBRRq7
vktpuGcYbxAZAjLRBo83T52aw+uR1Wvk8Z9AKWc1ZOUxql3ysz3CjWz5nJMOgo/wUknrftYGCk/I
zyIz4MvOGS03OtULk7HMOKnmHhrrUPR8wwSyU6P0q7tFR3QxPnRS/YTcvOUbNk6mdfqTn8RRpVUy
trNQ0qOQDQAH4S32KcAvnTuvlUVSEoXJTxupHv25V45u3HJzzQScwn2atqBFpA4eBHy7LA5Ccq8v
Imdy4h60sal8iR157b+g3kKeqgqskEJYZ9aKUUTsLahxF6uFZ28gqGtY91d1cnHbkARb4gC9YKGq
MEDNRUhubg0JJ9KRU2kpUT4GdtmLY/s2W6etc8vezKxiWjzVEJNc6c3bXhWRsGdLOoYWIfusJQx9
U3/2IkXxSlQnLvtvjuGTJDITRvLqoNgXe4KM9lkzJJaFic3tfIdKn06HdzpzsTI3YXzFeVAiekeE
hML+6WGXMVL8KK1rrXIIKn7sPv+DBQgq4WwImwsS9cY5ES1ZLlSnonaqgLP4n1ciQsUih92mZWXD
P59MWNOCaIm/FfAuJismSieW8L/Z67e++iSA3MjEOf8duYAJ5bLFDhk9rkIx252hpynBx8LEWrJO
I170f/5tD6w6+9ag4oi3ffZ6d+/FNeHIuweoXOf+K7cpiwBA6uryuDM+/sHAPMxRXS/LUNdf3CwU
JlAj6AZJSIoo3X3HDH7Dmhnvh5xn2nxK7wx1So54ksjp7vdB4aRIG54ZKvofrp9rlkoDRyyTx5I2
BeY2SLrdd4y1JvdEiO9tkjDePMwkxy9qqTZmocaMwkO9SXteGvmsWdBW1IHdDwKHD6zJmET15GcH
y7f08Hre/cmwizLc0uWzvl6dqs+pzSVEQSgIO2rlmlZOC+E4CDNz1M44QrADw5dGNFMkAdjz1L/9
Ssoy3PXneddefJcbVrYE49o5/p/k5f9IQjZkP6vdtAz+oq3nze9/gdVMP9gi+UyzIl5SYbbFbmH4
QLh64Xuzx/AFdW42lv5fyNwQO1QXA3K/dTjPIeAxHBJrkO2twZnQZPw+oquU83Va507SnVUJ5l7P
aB5WQgn3J+yu1a6LeeXc8NwuJ4oNgUko+DegEGv5dfoUdI/MtA6s7oaBVzYUg+0VIeQ3c5+3l0th
5iqKCpcQ6bBWSNbpCXi5A8RT+5jyusxFRc/CqN0Q4LpyA/8pOmAWGrgXJm31ABp0mzfgSh7/1PXk
meGCrhAsPBoR47bZrzWkvQvmpstu3UXgv3RDNhUztE0DwWuU9uqBDvZBllAMDFlo88on/D9RS0e9
efdhyJgqapkAAAm0pGGgD0l/r4a3287eoRiRwTpmO4Bw/L1fPwsDydhLtLrQNl/AQnHtrg/nGzKP
A1CbM+kkWvTaHpKnIs9jdxpX56K/38idYnVVps8GLDU7J42br3qgpu2ceHPz1Ka5bNIIqgpC9+1/
Yq/WxLKGWrDotGVdmfzBpkxu5+C4UgEtodNqxfMgwFSL2TM/mLIdi2rvp4MGQyIN1q23PqE8YPf1
Qms326ZiroKg9BGfw5GfwX0QSixtvSZZVK5mpkc0+X8W4mWq8QlZKH+r3DJrvOBu8FeWEGiXTqze
UQAQaj9/SPYXsEAzI3bunNXQAbnQpkQmsXaP8yHXN3/EwxIR4Endv+D9nfpRbTKYSCMnrWc5CASH
ySceuERBLQj+d+tqKCBsQ+kWrA7i0xflaHAE6BGcp7D8CjYhRrV/nwS0ssOapFOjBh+9Ca5bXTkw
xM8s/eXR3CQW3emZ7HoPjkXTtLN8aAIM2aeodNnqxfgBry3zOR06SlRjELmcgh2XbN55uGq8jNvM
ixVzBLp1IL8DMM7O+qzqh46etsA1zHbU+lZdOXBsKi+j+qk9RNlgSyin7Sjp3Q2RevBBB1Jtv+hW
bDO0vl7yScQKZNun8/18zjbOqdkZ+4V9UJcgvrL7NoeC9n6GLfkuP2AJiiKWArpDRQADrMcue7Ur
2EMe1ppR5gjUoZ+IhEiLGkziRvRF4YvaX2mLC6EL2JoiYYZNmnjygRFS+6ojC0SM0gsW900cU1TK
QIrsz8/kmNrS70UAm0neOA5JVzH1idaXEgYW7SNlmAVjTNS3EOtbNu1daE/i1A3pgua4YxpfBQ9c
TkokPqixy2wsR3RdWBH0q8yCEMTfaekspRvDDbwCea2AL79EQJyDf2+luZ5HLQtNGozkceuJ3LJU
zY3N62GESC04LuRwbtfrd6ydZvnQqE6yQzG71n1wbwccWBD4lTluAA9ffJZobtV4Qo7u0rFOL3zB
3Q3hZDXPIbEyoQHes4OZyUZuOoQJY3BPyWcza3D9Y65hLt8S9aGPy6OVo2JS9KAOs36YtBoKLH0O
FiPrXlpfq3PJq4E4vuKNp2CVdoNLbuirh0oomNhhhvuFF0hnssdSgNUvkvR5YsqNLjtvuQK9KWnj
jhdRc0FfiMJFj9xH9Sm7cU/5ixCobkwZYYFJn+WWG1qEcNr3/Ozl97DsiWgbwCU6nGxr+VhS0W7/
zcUeVXPxY3/j2mR7gfjM/VYEhMpw//hw506qilPdASAZH+ccXrogxXULR4U0+iblH6dBXRvRFYgb
YZUy4GnVBrfGBsFuLoM3/9YEsqGbOYpLozt4L+ymCZ3nH3MLdx5c+LEBix/go8OvJeTmV5ki3wJM
Xnntptm8KZCviicIrApBAr8V76BCarOdIyDA76HynlBx00pYHh0kp1ZPMhRsBR1Zh9nRgrewZexK
u+3zlU5w749/mCAc/YCLrdHz4tyYrD/sXI2gYRCXd0jDxDsvtiKhfrG4Q+/4UgjUGzVEfhDUBPGN
rRGkgwkxmzLLCNseZAnqTV0yUh4Ku+AqSje80pXqdd0tXC049f7Jwr+59XpaAF+TgYfsIep18v5G
gMnEldMMKJUMJPSkUX0JJjOxBXcdY+cOwbLM8s39bSPp9Kj3ip+Qq/r/pg7J8nUYR+8mq5BfA2M4
o+3nwbfmaMCHf9Nt/jaxtXG/xPqTwPtfGKzm7/o3Z35wVKkGF+JzqfwutO1okhBQeCMlU+TBGwKP
8SY8/ZqpJ86rPbbsu0jG7mcH8rGELIP6ch/d3TyzdK8Zy4fe0oaZncy9xMcRkZH5bcqgLmL1gcMa
OHWX+3DAqLkxYiShsyGIo2uN12+E7JRZ2TwxS1o6R3O4iIgXiusnShopZrVLwEmkirqwosAyNtNX
ErwitM/Ycls+OVDd7Nm04CcicTjJoB2ebb1WcBrSvBj7iyeR9UBZ2OWcc0MXvnT4dFfHiPV7fPtF
yVqYfRwWv0mAWUbcBrhu+tg0Z/eL4hMLTMZmaHeJ93C6PDnos5sZjODCOZqrFW+YCyezoZU9zPBo
yXwBU3Tq9QlSIVjPScATSftfFkZfbIRaSqmTxMza1luqr9rbFklVwkeEGmCy0xZf04OMmdshlAXz
hdTrmIOXTzSp0gBH1/MVmk5dT/bAb15OyFn20mzeuIurV9CBLw3B5Xs1nH/5MuGPQUBkUvAI3gcb
kZI0xaAoBoPQh18PnLUkzrVI1MIpLukRcv+w4qElses5fquCPeuvBmo5zO8nRHNuHMwlNcsLtLXd
4MeTaljYBloeBAnpXQtHB7nA+w0Gi8Xb/ch+kpa94si7drijfm7AARmI9bA4ZyJD1OOI9aEE9qf/
rnm3QtHanL0dl3XrGytSSgM8v3mmkQMhzA3VTdycndy06H5Bmv2q+a8xON28gELJHrLKk0iI2cNM
GMgnTLJeYmRFMPQEWEg5vebaI8ENvEjS8P+ZA2LkfctiRJADqKYmKV4Qxe1U/8mDISp2ZKA3PEON
erLBhKP261YXewhoOYbcM9KDBTWq0JR7EphLif9KX79OJuNVhgLxR33OVfX9PVXyxMptSTv+boMm
FZW3lrjwOldVrY9jcpdOfFEU6GqrJGSBhfn58yh1xVsILoIlr8tlD+5EX2BXnr/8Hr9AydZuCUl+
9V3T46vCjNj2g4j82YNHnnLDjok/4J2ma0tM34Q83SpWi9Xz3xcT3mkLzsqnQZ9TNfzRp29YNXsR
hLep6FxeYCMAdZUGpnAwUYQVg1mZ0hdG6/gd6xXQpJR9/zvXPWlinsEWqXkUcri4XxZS4yIcCtmP
aLiooB4U7V7PS5TNoscEsdoMGbqK9Wc9RcO1FyG/0/4EzAbH4sFOM88scpVVDEoYlXsDebEdfDts
sqcX5eKzTNMEmgYFJmIhtsN8dhEuMvSBZdzpy6ygm+v2Bhgihapw16+lp+Pg4pEHQp6LFoicTHN9
amxBiErTVUpXXaBXDdG6MUhVc3HpG5csLDARMhJOZlvJc3FCx0zriYonNYhrlHzzt4RAfS+38Jcg
9tK4111HbmnDVS5HULAVnl+OswS8JcK8TLafeSzg63aCT/exWwwTV6uidYBq46Hlmla4byDr/UGW
VA5WluQyImRMS1rkNZ/pQKkw7qU+C1+tmNXLr0liXCETlIV4DF2DPbqbehLN7N4t4KdTc+9s9Ish
ECjeaRwtzuZ2TgMpLJURS/d6lP+Iy1gJWcLho+0mJlrCsROtye1bzFVCbGYerB89nk2ejTSiimjV
N5mlAqecvPkdi1bMdG3h0KoaOlwvQlfDObge+Y68f4fSdamVpATfnBTv3UHN+oghjX1/NAiAgWp2
++65L1KqCJmpALzS0smnVxQaXFbIWrFHn5THYGuhgVhkf+9CSKep2VKIjG2MfmdMvFj9v5HdRaWT
pcy/LqrL0Fb0KbqRQk5UGZNPnSiIZHXQHcTO1MZTm3YxQauvxKxPlxs09trjJbmlol/fhiCxE0DN
hqm8SfiDxvDqPl5ecAnsGLw1HJbJ/MY0H527/Yx8dM9PNFBFGrX1/0sfqp26X1BpHVOxw6iktp9V
sdwWK3kHUEwqiv7OhtmzJy1zYYaje//+0PfPW+MEr3qjwKTSck53BiGyE41J0/5YClhNGtfSjl6E
G4E06VS6vl81RNB/24BwBLiGTn7Hy4NTL+uCdqoqSIieOBMaDhsK19gefI9acOxdoaEk5NkCwBck
edFC6PWtykh5EOKFW5YKG9X3AiyJ9oql8SAOXOZvwNsAa4wZEFCf54Ng+5h7Izd6QQ5RIqJIWS4U
uzK0fWIRkLd7781ZikI2gc5lNylFVyic+kFnOQadeJWq76LGl/OKlexj6OR0z7qtC2ovNUxdWAzg
/9Skz2ZiGZvrWqus+isQuIrmc2B3cfiwu6ZPJ9UuLNTAW4WFeWhmHLQzv0gXHQBC/V9bYnB8/kfH
fOS3OO+mqTH1KKXGCiWyYGpGh/syH2OVYjien7NxsBHR9NG7cbihOaalWxSVATQgFxJq00Jqq9Rf
OgWkyNiSDV/xtCSmx4mxJunNk7zmljEqfM/pH3zMWu4/6NFNfOZA4X9y+/ABs/5DeACD6gkuT3hj
RgbRZj743jG0TwZpHcd5o3Js+25tWRS5LDy6X10G5qRfP5y+rsrzbMmhgSsbfRWVXw9u/brYUmcZ
sjfu7rBi2OBD9qiYherR2lj+KnsCAts25qGwoCCXD4jqx1f/IaciKM5BRiJ5lhBRFzaHpoy12/mR
DXZBcTSY2DwRCz1yqeo6fulhbB5GpMUzLi7gtZRbWMYUfeR1lWcxeDcYdWYL4i6HhVzUfTqJ6ywX
QFeIwbEF2HgwJkeloyeeEkqvVAc9jSGSoBF7EIOK9XmIowcxgBhSnLxDCRDTxoPrEcYshca6G0N+
7KTGfLyBqtRt08YFEG3qo2Gg0yc/I6BbAnDU9pS97pmiCQVK+ctETKoJ307cdpn9W2OsMIaVwB0+
ANexPKoJzcxIJiKrYlbLFHuNOsPMJ+XjK/wwowRxgrqBMd204y15YjkkgaiCoJ9YjT9vH0MI1tnF
UOeYOqR4C4SUPQNxOAh2u+sBhj9g6m8omrlDqlEB0F2DP7tmp0DFsEOmLmkcqcPGouoJmmyQ4UxF
wvfgWx39LFnrTWagAj3Vtk2oQtwYacTHieDCp3z+7Zycz/ohQQ9/2Vm+N+KYtatrQinHrjuzbWNp
I5Yc2TkIhXLX9+MEGmDOsu7Ei27Lzhls3ceGVzSAhmZlFXOCL89jSNXGaMHa5Fj9QeYW/cCuQg41
GfzmOXiIBL05ZBG3ViyhH40Kqo2z0z0qtsSLO91GMQanlIFLnQZ67tJTF09U2rLD06i/8DwLNFWr
hvbjvxmRUXlwLDyhXuGDpua9/pvqeMX4X9jt/wYbuQsDyUI82yyqnVmfe/8KyUXOhpdl3SJx0IYG
vPwfQGUFTh0UX582TUT7Z+PyP4scKrec9ImAUfbE9xeIP+wETBsBL9oXxW617GZfYzxH0CUIQHz1
v/0YjHupGUnZwM82VLw2ziIUaMtiDbZDzPU/TMRFxrqHTrx1xhobHIBB6F4/HoNNyEo4sejf4yfO
2n2OBIbla1x/mwDst3iRUWhRnd+krXPuTCkN1ImRuVD0A6feIKFubMK8vTddLA+eCHcLmKCJpHsF
T16ZJqj1FdYZy//I+Rl2gIG+USi9jqrgzEsSYZ4NpGJbwNR+isYJbsvuLkIyA84LEhPCFgUQA0ro
UWFxUnJAKC0/cgmcWJY6c5JAQYUmtzNwASaF+i/qng+n3RN7/VRcyR36P7dbQFcOKdsLUpgC/7Jt
bUbxdu/LR94UmvhYzSb/VYGLtyXK6aYgY3tEeuujTthji5vEoZC3Fq48DhL/hwfMS/5FFlk7JixG
LqnjxyVRO9fn05BhaiuNvs2O/6/ICChYZW7+qABFoaJ2NL6hZrEzOLvNO1oaoTGvzF2nhCvbBKdg
G51DsZajrV6ogSUf5RbHC9HOZdjV6IkakiohIaUsca5bjYK+CL9AgH0UAFFIL+M/wcW6JVqiWdo4
eyRnxNzFeS6qigZfDV0bgwRqmB+sui7iT/KFtsLvWoa5Vkpki7oAlC3tIGi1zGFcHQBt9IqBvnET
AUVRMfTL/rq/H8hVU332bOZbRFvnGjF4ryLvLFGdTB5cnCdJMxZ4a1sL3axrnwr1pnBvcKWPCjnG
kAAb7pCfB5oPxTABjf0YTXCwFOf4lvYmNK474xTssr6cvsKKBeUO537ycH/FYYC60JLybE9OzCq7
wstC9AkpGfjgN/UzlQnE5SpXF3uY/NK1LE/B/HoRFwmaZYKC7t/syWgzV+07Wwpzb5UlX5hJb54i
WfOnuW7lnMVG8Ej3weKnl58AuY6eo2R9udQ+qA4bAWEIruO5KCy9ijBFxg3d9OLhpgmXN3yzERm9
6q8f4pFpTcvKViSSXC+fB0oWTg1OShYv1CCxVfmdML7rHwanXAsUGJnm5VymJi7rZ9dSlGe7SbYg
ac92Pge1pbSQpoyP0e6gO2fZMU7deXcD2o1JItk9mj93CLGV0ioa43j4YyGKIbsR4+8GLcvevHpX
sH8Vxg/XM0o4lh8w1692tunoyj/MpDvC9+E7gEoC+FAF683KlVexMcGFKZhhqPd+5wVY35nPeRSH
hGeCf1ykK8t6fYnzDZXE/lzQYDvHl8hXMoRu0clwhl3B2zdUIyfhbmFUKBNzmRE6Hbp6q1I+H3rA
wJSJyTvoI5f1Mz4IiQeYqTpznTJFMCVWC8D+IU6KYgJqiZyU/x+Cy/M6ORWugApxmUphGSCvagLJ
6aEd/9FaCnt3Q1j+8P0n266LeCI9KN6ObtlQBkMDYPK/A8hP6oh3UB7ag5vsRn1RAcWOSeuyaLJ2
X1lE7K1VPYSvxQUfogXecuxCSm7dDC2yAPqkA/evGDVZ9he3UZ9htLpjh2pryyxtDE1XoGUkh9jb
1IQo0YFMjJLoBRoGnCaujMwhGcH/zbMlfcfbQy/QEd5ICRzLsE+cCKcNU8ddgYXX4rn0pM6Lx52M
VT9tZ5VdV8yErPXAVYwnk7mpoOsUS8u3XZa8cCoQ1IQbfIrcHKUdT56VZeVO3KKKB0MubN9SAv4M
khUYrUHnOg+EyU64lgY9e24SDyNGIyY7DIyNuglxntzhueSvKI2qAnycWRIWEn64Q/vTeOQdTBSy
lanFHvZxDXD5h7bTiJSWETgdjotZAJTfbyheSXIMk++xWBi/cfUKKjo7/TuF7XKVEFNSWHgsYeif
xPcodYS5krMzM8Sz4E6u+1rW9oNXrT6Ah+xCIRtjPTKfyPYqTJQrgJGb/Vjm//YGtZCx7E05/dYF
sVcSIyQUrMST2VbKw7oRmVfO6yZdooHey4f8aBYUmDMo90j2x/7AtKW3punkg6rADAZQ/mgG0nOk
b8MGcd/QRTZYFNWHogh3bIpTzV21g/J46w11Y0EowRv3hCbiPAEyJWnNgaxUadOj1rXDbvT9DNdy
GrjqIpBxDFVz3xjd7IID6ncctA4eLJ9OFuRm9UVyOFVGuwxCULAXaAayijV1+NrUA2vuuljI6bsf
pPKTQInGxH2t9JcTf3IYgXJbhaHJfWrw8UiLtz9E4oqTe1k7eShqtiys15K1tqZz9HyG+cCZcE98
n7hWduuqp14gR0Gc93H4RNy7o89tVf7ce85L1zLZFmOXSctXjeF81GiiBA5MxTQx3ZpLjXpYQxKO
KXonw8LZtg3UePN6guys0+k0fhRmWsWoCVcuQKlBwdNKIHUKyXeFX+/SpcYTNjmC8/5I739np3dG
EshOjRGkc9ZGFMtlDP5aOBGuRy3EtdE7Nyefm54nGgIwlQ8el7gbKUWGER8ZYHFmexFk8neJV7xz
jqahfquLgYTR+Mm+ot6i6DDLI7RzY+QvrcIsJTKrbL1N0I9TDwmUYThHYh/U/zS1+jHoe5Fp4n7y
RZ4uoqs2WK9wuA3mBEYcbws9t41HrAxTlrKBSQZ72saQxFYRiFOTvMh3lEN+vEwWoHCAs3AqD3RI
pW4inAk8TwHuGRQtHxcMdroyKXDCoQVry5qRgYDCWtG+u9irIWMgB0s7GlcmKuC+j3FeCeDEoQ1Q
04dlDQclrD+av4gNdYMmRo6Vu76kuGxUwcPJERJEIYVQ8irlM7etM6zopHVkDnc0B4pMcrcTVLz9
ujax1M+yMhO4qPWGmFxFpCTjESru4o0B47PwKwMq/zPkC5CRbIiJMByjYk6nNuCl5zfnLGVFpN1W
5REdcLzus6jyNwkfbWEKM72UZC66L8GGOACbnNP09MQSOQLM/tnSoCqBilDRLjn/+sRb61MKoMxI
+dlISu74IEYYFrJsfOppxiAXFBnG4pU9TYOkUb0SqLLhsLvU4xD44wx8rEtxVQCOXFgolv/6I1xc
wnIsuy9OJyEMpbxhPO+n+5/O1yYjjpiDiGXvHL/0R40B08wSSJALYVNdMxlzgAn27Dk1s4Rg9zU2
q2yURD4SQ5j/egA5qtAtX2b/+1cYQ9OYy7yhBdKm90wJf4u1wE39Q+rKXcyD1KojHc0355ChKKis
LAzfAvPIDSJBNS3vbX4HcPu/CX8D551Rx3TpJ2AwB9FFX2wNKLNM/eUxy0wYpzlMBYZeMn26gucD
1P+cE7jChEZIz7sBSogx9sgHJ/OJXRSsW0q4jCyHW6E1N0s/hTF4R+GuVq5g/Ezw2oW56KcRNM6d
psAajnxmSE8ryK/RtE8KA7aFYFYNAACDcdz2oZkBAYANhYIZ/SG3V6uOxHWTUstyIjp3y7yoSAO9
fOMXICXg/WSpO2GOacbO/vGHoTkT1dWjF/ogB4JWjXYVH69oB1yxSH/MMikLMrwtZck1dQq66nYq
vQPE11yqxkgP7xU48MDlYP253i5Mqg8SrkFIS0bk3GntfacxLROoBey5KbaGZzsHUNMgmWQA1Zf8
bhVMta5Pz86uQ0yXSRrfHxFpgPSJoFPqoY801NkINNKYRD1P8MQ1Gg/UqM3zckYWnKXNe/iVkVy8
MQwUETfZ64HvHnFw7EBu/+COnw+jMRDzU4nANYK39pY6I3hQCqYuX7JtUEpBL+z9gbwHcqPvwnXA
ajvZV3cMnhmIJeM7EN/v+QeFfmwL7v+NwYJ0thv5IiuCwcUyppBSFUaylpic1G31JVnApCVycuk9
qfoFFxDgRC1R8c3ClkoKimLD6l2231YqoHRcobh1WLgKqgHwpRhgl90yoc2wN9jUoftjD0Vp4/fA
tfVc8Ge8cEjcfGJOqkxmzcPcdOQZzHW+qqj4lt+O3tQ5AqXDIs+rUaAjFqYVAHWUjwpJAhPUwKAf
OB7e+0GcfoBA1KMUQRibaqd6afei0zLnMNSnGbX4Imaa4jas6hjsw/VbIj1zqOG2qpnPP1KUyv5F
rxLxWsYtn0r4CGaGvqgD13OYzz4B2CaO/defOWtnLVnZBdBVg8SCXM3dbU24jgmbOm93Y9McMuUX
d1100/xZTSZysptqfG5zIc7QHHDZjw0ixN3hUaBHf7k/J9GNgVAlKh3rtPyXJnkTjsuyx9vBTwEJ
PV3SVG5f6o3lEcnnW9oREnuL328H5rU0VckIfUHzC+8zPQjsLIzpM3VmU7xRJjx1uf4ERkQ6kU49
ZrUI2FHj4CsYCtXjZtzEqQJ5Y4hPXsp4V3Zd4hRj8EZmhsMXbKEgFzOnSDTWZdQd3duU4S03WLZF
nBnhkSbGTw4fCYvqyPAYTw9+jKRRGWHNV68fpsZeeARfhhytiJMfs/pXwTecP3FA9RjbKLeSyMW9
AcsBjMKk4OxKwsiC9CrCT0PS99aKv945wzoYNo5J39jWgHIXPavWLaom+l0NlNiQtuAA402llMkL
RNI4qSNbq/8FBheY+xhEaMFNBSPRVCTvaHOvJcCNFdhNVspehRwR4yxiM6UZHsfJIUPaErnoCYzu
FJqprXBVipUY6g2Bjr8V0DJ3FVK7xGF8A/Icag/2uRJvKTInxB0JS+PNaXd09ensnhypUKXLh3w0
bJsjp4PxKeSBTxouPSFI/gJhD0irMUmQubG5RAnp+cG9OxEsKvxb22Bd5h9of1NOkAYsox/egqHw
vdiyGwdr2eMpUdfcChz6QavNTG4NBJpflVMLYbPbI2Xnd0glYEJBj8mgXzKZMbwTePHCPK5ICqiM
2vWw06p74YSPsEwb8C67MtSad6aY1WdfIkLZ38fHwFYdYLP/YGjnfXAumGM+157NKpcFAD5P4FPN
QvJw88EB2iNJ/XukPMLuNpvBM2kMK05wS+SaxiP4I3zX86R04JHd7ATYzY9DaLftbHOgv0G2cPfp
T7VvOESAXth5luQbQPTP8Ko70CGSQ6ZtjyVkS8Zhkfw2K6YRlP7Dv/QTtAjoc/vzoi0JrnEaxpPD
wGtUcDTHNnRdxc2Gq+x7Pr4cm91vYbtpQtsqekFuk7JMBxRygor3p18xR5+Pk/+uRT4Qa/pkSWBx
i7dQv5zG1IDfspmRCAIcoPBuDJARryEUcoH4Th6sg1eKAiLNHPZp0uhGC/+0FXac9z6YTovtR3Ov
O5HsICYP9SH/ETHtdfCF6h/p4nn4eLJPCW7b4y/ichSvBNFLOF2EUWcgK5iSGyC5txaj8S/1ibCF
gg3r2y8eJ87InSBuD6BL2tmg2r0toPGd3knW8YKkOG6q2cgcb8qqeooXl/cS/N1S2Z8K1MiGcghR
Dl622d6UHPRA8QHHl6Fcwwm2AICl00ixpjUZq+8VOnNowRIr5SNm8kEsLqkCDAeygjWQRT5ASgLk
h2D2TY8xIjXy/Mv46xC159GJcXuvQNN7wpNH+ZxbQwZwNgSFHmkDPTCCIIzMmlOxXM2t90HCo7QH
6E+lNx46o75tCGMfGDVaToZPlmDEn1i5xfWBivvZ99KANfXdJK5H8O0jvf9HYXKE/arTwm4BT72P
OfohpgI7V+35iHEJS903T1evcOFvherQLesvwPvdBUqKdRNtuEKgQ3gcj0J6tEAtCvgXYmuCIm30
wTXjKH7qI5ljYT9rCwLHE7valI667RevlbW1V0lJUx3Ugn5QKLjc4GDFgav8uC4vbb1AxESwJyFI
uU4lt3KwD1gD6jTDYtA4BIx9KEorP+lteuNenLHJonvbuIPF/N/l7bZZRgsHuyOIx2bQPslUi5oA
/TBB2JhRQz0fyAu0cUli4j+3gGAXygD/hp1a1UuC8/pdxGHDB9BiuKtSjcoDwBwsCrajnhb/wGOj
TUmsS9NPW6wI1/1Vwe8MyCPHJ1REni6EuBUm31pVc6WbRXMu3Rjy9f9mbsfJTLqIIXS+HaadUkVK
+ZXWnvcFmSM2/+VsupdZn36Qh170PH2uAJV3E9fNxEpJnc7KSh5Io22lq3t41jrcZr1f3TTMMAeU
VQJDOZlzM0NYuZ4MJnpttFicRl1RzTpG6fkBNB0IQouO+bPSzwFTMbbSHKEeDYN3ztjHXaZpIbE6
Ro/vJ9Ra3sfdqlvz0fnVpSd1rUvhwgY9LmeLRRsVWx0BS8jqBJsAPYbxHMD77IyuUTCAraS3dM/h
USjhOc69/Nqkl8hvASe3NSyXNh5R7boN/OqGyMHQ+9yD40asnTPebL8QAZz2+xNEyL1kwFZ3b6o2
1vRTqIGbS5UL5ymDM9SDlcjwfKPznTKhZ9arkTzkgbeP2AlwM/ySODIyKmYzNxg2LQSmuo3dWDdG
7xjtEuowVgVZfiugMrvf1MgD25SJKPcviWKNSsgi+ffz8NULWS0jiY5OCZZh004S1qPgWBEKzIsZ
HyzC69medQeHFrIa+eHrK4Fevwza1wgVukZycAY218/tuYQ2aCZdKQUePoefqVgcRr4Tn9JXj0qy
23EFeQzERGdTj49LJYhYexi9uTSJhB2DARqXX4o7LJJ6uyujTK+qHPEHGz2piqZ2qEDknlLLmGVY
as5/OQvPkDHIkj6wtik5Fg1to6npzHcdk1BANea5ILlSV1Rk9/aLZfp9a1whE9Hqu4GFsx2UYRCT
eWSdXsNZw85Q6QHdq0CLSJ+D8UpnB8x7yHQo5+vs+v5xB28zuWweD1Acvxo8RqlcSPcGg4JQ6ohi
q7vWdwV2fHs8g6JhX3RfajU8NbWTbHvu6dWaEfV3+BWc/DvvMfP9q0a07JrtmiUxPmXvIIxhX50w
0ImiMLIJHIwmNB8jGgxY8Z7WpABpPZ14ZJzUQvOe5SIR26DXBiaTJp6P04TeDkP4EP7wjK7X63EO
aWQzLGgrbkHcO4GVhcF0zVvfuMKn7YJj7xLUqZsmJYpRxQC95WRKNzTTTTU6nwOKdiHx5aoOJRad
xljCMevnoDw2okkC/7XIQWIzQN87g+Q93g47y6VBlHGOcZZUMydwWfPLwa0Pk3jM54qrxZKqmBjB
dmfJEOlahxY71zHpCYv/7JoTXjME8kaRnfwuo5wiIpFZlV3PHix6ERtSk3TmWc6sjgva2+UiV6uL
kungXoFYHnhIS6BRG4P9PxWbzs3EobktNPsmwGukQi8/hXtksv44oBVNqsumA3ir414uIRwt+K5u
dUMjCLvVzqIHfBXAuFpYtaR8xjp2zPaL/NxJ32bzXXmssM+VFQsA+LCzval77F1Z6oxPYLWhNGS1
GWTdskT09LmF4PUZumcPyF1EO1v/Iv41OtA/SSeBNUJQqnVj3IHNTMB5yP2fVU2KiFMdvz5MaUc2
dIu3YrGfgfDQbdFz1SNarsu3xxN2hYAMVRV7py5DwEpZSwchSWHnnZvEzsO5UvUj/b+PSlh7dGXK
bhQfg22jsZEZHAKus9ZKrr4cFyRaEUOKU3Oh+099EFCr3zivb2OGbIeIhcyb7+8Rd+K000zyVLGX
GvlChQOT9bcizfxJqeX2lxFazLs9zaIUCyXbCNosynWgRbgejjSAoTygcNvPFc7hGpzrewN9GqYf
5PSI7ttxWgDydPz6S8qfnx2yB6tsU0xefQqvOpzSeCCPuSviuoUq1ggveZjitgPxMFnSJ774deNJ
GkiIsc7FaxddC4EjUlAdhmHEszs+nCmuO2jsFwOh8eC4e7K0QT0Ve+WwR2GefiXMve+TNyweyntj
NyNcWBOVktcXuQxBX4L4cVvouaIsJQ/epQDB3QgFd0Ty0zxwIm/FzxIF8z2NbjLFIBbp4mEXVahi
rYsIKvKY6tMpoRGvg1DBvsg/LoynwsHUO2aqZwPa/M1GR9x55kUoiX7R7jGNTY0u0tnVgY/iBfOX
D0LpVvdr4H90vTlTfqHNywCPDKqp/Y3t84npWm1/CfJVdttS1C7XcOjHrxyBZYHG6PZnoDaL2GSM
MYIoPzHJMLISIWqMm38++Q18QVeSOSZcDIXcOEduQ2h/AvSyvUJVGDGB6EpWRaObnB8/SUrDZUdr
k9E0QaESPS7tGAqe6Njx/l6hdwIcuWTpvvQqeBLNIVb5YPtg8Zs6eHmk/9zsN+JemhtziB6W1Ykv
mw2jmcOqeH/VvyM42M9nXEXigPJm8z4I34WVSb/iOw8qQFRjfe5ZIrAxpaDwubGnQtJMtyg+BfnY
OQygCmPJI+82Ehr1bCcJ7cQk5gY17H+DxKVqPp2S8Zneb/pQA4ckVHWIbILBqE5Dgewspv75KET1
a8w8yWPCmosn0NY48c7r/1tFG2mpHeUZjuSZxVp5ra39SqqjeqUwxDbLLnbXuMLLW+/YuL/t2XT0
hVvfKygIyr1QDOF/CmQbEAUl2OUvheu6DZmCRdZl0GcwcgxAzIDT/z4RUhoMhiHY8sm+PuHk77fI
mSz/kA6lHaVf4WcBEkB1b1gOKY5KKomL7Ix3kJYdz7PkhTI6xDUmxjnHYfLbYxTNKrYf/fNhR1RF
VvqL9cobLNY1bhoTS6cAOJK5sR26retUkB05Bl27C5Hv65XBw3vKDpwZiMaS3Id4OCgO+qQLjXWQ
a6vf8a2+1U2tr780ImQ3CoQKj0+hF3Rp/NWiDZ5eJot+J4O40uUjlqX+mY9nXyPJyhrRd8DnEc92
dibXyuU8qmzWcaxuLBuzoTcAhmTe6XHfic+fGxRcehL7xLMCkPkFjv+ON19wzoaInlYRUsrf99vq
b8FdW6Re1Ipi0o/gMj1M6e+aJ/Aql3EcFq1uPzt/pWwhjRdCaXhd2kQbBdNA5StsQiQy5bs5s4M8
J4Y+ycqUylxlJ+9ehG8bBMP6VltN8AW+Kqh7AFWw/ADGsBezP3SWeQIXySVHI9y4yykXix3SA2yf
VFhnnQ8FlnJe0XsimSDGZOcFeInPDj9M6YyK10bQOWjZm5ToRhNohYErSEzJUMYlgVL9VY2Y5lkq
yNqgozDWxkOGXyk5OzggdxiO3xwDKLEgTUKOyf/YpgZAph8DrEnGD8TJtB1puGScNNa47q+MRwgJ
Mnh6ot3hnbR5OMslW3bolZx+JCNWzNbvtbJCHtlXVO2559lcphlAP0ed3+LPVODq1McnIzBs/Rtl
HemRogd5dlmHTawRlQuxw/HOd80snJQoPtSfBAWvxcHHmQGMzYQRSnesgoNj3qqwJQPQRKHEAobI
DD5xiGKR3vYzbKBKToyajqemhjXO+EWF+/xPLew6GSXFyuUbtwWlQDVUjh0qvxOlmjlkr80haMXa
lLcpEh7CML2S89friTEeBGx4Irpcj+lCwgv6qkHSfPlwd+ZzYusWMfDU4rSKz5QeDvlfW6RAyqL1
vMxs/XViAIROSgpbbrF00/59pwTVr+q+/kotOhCsW4Eo2ZdaDOiOPCqZpWLXInnvNRhTadqC47b3
AmYo3ZdxR66Rjrm+DRIVyHG9mFEwUPu6YBlRfe5+9P3X2Wk4ZJYv/c+NjVSm0WCtuewz9CuNi1Zy
rrKZq2PucxeN6SNRjcx0zlt1HYJbzyfZZS1llnZ3dGhAlzz4eOZXX/aPgm7K5o2z3UkskNBcKwRs
KsYJNNeqarcquJ/RUMxDwWiSLhUDBPa9z2lX2WIeKPrdWzY0tO0FFq01aFTZg8OAtDl/8wzDyG8x
boiqyCde6kIfU+VuCrrL5O/Oq1q9ak4BgzK99VYExE4p0BLdPfbvJwS+1n++PpM18eejBWllrAad
6M9S3nbzHWipHbCnOqKWXjI3mqpPF8GaE9HsyJKvU1C8ae8Jif9dGk/dXqRmTkyYUfjYDQPMpMr5
Ii88lVH+1HO7hDTNWMcWw3CZVUxTyrIulXMHGotPicXXQnReOJC2QoFhsQwZ8qFh9cT170mHCp1X
NWT4bcBkRxZsWO9CmNv1O9bYxKFPPa/xctSa8wAYVFcBHDjzQbD4N5dKVjdIPOgt/OKaQPlMk0NN
CW6PBgYs91uaq9M591ykjHTbuTYW8BQAVXFp7MrqT0uB0M8gmPFudthzYW327OWL7KdAP130HPv/
70S1X4GA0BZQGaawCKvDSxVRwfGkpNz5WH5kEK6lX4TDtWbQ0cBf70Nlj8jQKdGEZO3naLe9naVb
YkxNYSw9OykqGRmze3sqG+REJ8DVmpkBYGksi69Wb+jOZpNwfp1hVmNvMtyjF/xgHH+dh4cWgR/l
+epeK8lFPHgN75NQ/m90rZnAC4iUH5epICpnrjvMGjqx+GJKsO31bEC03vJgyq3DXA2VlVB/XqTi
V9PH0YEf5kli1eiNINyXKRIOLrgjNG1h3ANvAoGB4CLnGayms4xHFi18qZfVi5s/CssZAQ5FtsNM
K1Ons0Q97qnNYUU1vAYep++nfkMfAMqFME2JrEpc7URexwuT8r4uYSxKoYjGLjshmqXnpRiGbCie
nw8Tz79OoryC4viWVjqaEGiYmUAdpAy9E8wvV60dG1iAtZgtgngMEQ2KLuLz5CmMrLeDWcIxWJlt
59HW6ROgLg4i4fUrHdpznP6sDGJFQXylUEpeUQMEYxZ5lBX9wNHguppsb771qb+Jiu+MLzKt4Bv9
p+HoWRpTtHZtC76W1b/I+A8BUWDQHwQ9n/U2r6TDr+65WOz2R+6WuUIVXIZJnuo+P3ugjZkHSYDA
K43xkzT1kLLf+spBULiFqzLcwhM9UCH/J17DUesJbOH8tuu9258HOcY7zC500A3uFzzUnWO4svFd
Z+e+Pv+JSlxROV5/TH83P0Nai3DMX2m2NHqrXjGKVPcQQ88ZFNACwVuATv9acT/mpGYH+1Q14xEe
Nk36/UneS0xF+lOVpERyClFc8uIQXVcwCEfRcwXkfdaIbRua7SMDZcpgpVBlCId1R4HNETxjcN0m
AUjp+mDyR0b36u5vQMFnr7FKJOtdmbKBRI0dvg/LmYeL9Ag7qlQjpJW4LruXFv2PCt8thcJAlITs
rxYzOznAgGM8RqOYNLxGUkaQg0jNf516j1qV9GYVJtSJRX/xn5POZt59tMSYbcmNGUYvyuXbV6k/
KrRXkQY+fcoz3HH0a2WOwQzGuOfChfM9nkJS+5fhdiZ4A5/E1Wl9tahETPzC5V/Z2DiAl+oFoD/Y
3FeKXUvG6s0ql9b8KXcOsUebcuidjJWbe5VvJxoLFi9+ZGJ9ZRjZGbds0SaEDWrowbUpQtgwjJr8
vf/hm7EiiQzXeVaF/KMV17vO3pCU2DgmFOPwRZW6VIINkEMT3u4cY3BqJ8LGINNf4D2uk/vMn4W8
x5eTKcol4iKByAhZsyae4fMvfjTS2SANy5m5TvAWBiV6Ct9DJm7ZxSCpW2kMyPtnKo61wYZLUTd3
gaaI4jZXyUQIvtTo4UD3FHzVInkOdoRO6LJ/p2uJL6RD9qIxv7/gdw0DZ/lR63tvcuTcsAp1u/w3
0Gu2DoYaJSGRz8KUSg6NO/BiouUvDrxLiR6RZpQyFQtMSCAKPpusw4n8uEB5SWYeKUHofwYJujU5
EJHlmu95Y5zTWWtnU3dSsftsv1bOdqEUJkHOaxVMraviWksaPQy7vRg9jOsCEx5b4fXXCiT4xJx0
XUweu0GLSIucAnw0wDKuXmLwIFSVI2lQC/8Kw2G17CMKeD2c950bHhTbrLWOuCD9F1w5AHTApWW5
vsW4kHFj6qIaoiS8lpR4t1FCttYe+B3HmRnzhnZlEcHQTPAFSa3k0DNTLGoGjhL69o4Ol+dHIYld
zolOWXGcH0o/IhZygL+qdiLskYnqqXTTQKdcQEJquSe9VDDAZoVe+bAXR2RAzDW1oPmnFBgctUd9
SUkBHj+h5yZxV7bIh84DKJ23XS/7t8y6iIpVaBcPuzUGxjRIESnoDq2eZn2Mb8HGUJfGy4MXAtzp
NjxWvHgQ3HVD2Ct6VDlfBtuOzprhdXDnUDc/LJvvVEArXImF0pwH+NxZdU6gUQMTHMpOoxfOCowg
qrq1+gfsWRFMqeBhgyEzsNak23dP+Dt/WAbOFASFBE5BDt2ZChQAKzC4zo1Qsa7JviPTqQJp515x
77OFc0nl8Pwo8g6fvlG94yxhKzOG/ox2sc9YSDVbKETgBRtOnYGrRQ80IKOCxP63hhlMMMtO78pc
6EvrF2liktLYQp8hYCwVQYJJc+2mF0rjNkVVpfL7Pbi0MQNse97+u8KwP01j7owRSUKiTu+WegTV
r+ALspfO0sspRyl110Ith3S55244eZ0N4eaC79GaaPQgb/toXg2zVFrl9Js2t5UxBuhSDl9GRN10
MCwodJ4JlcQN+bQOh9eWnb8uUIbaT08gVNIHXOLOHQfpX6JxlQMu7vD6N1r9NVWNr/vXgyUjIFKF
eo50Q9MlSHvUqUX5dEUdkz8bRgLIWU2hS8ILdSBe5KSEnkBCsmvlY4IwGCl0LwEOfBCrwd/RH0Z8
WtShcw3tY0bvuiHs8OkrXusyZEm11qIJqRkFcQmN6WPWFy6u7uhqxzZK+FiLJYTQ7ccxf+ufB1k/
JQZtl6Rd24eXIoKSgWsbJLTLZ0jNweNVeIH8gfZeMNpeqeihBLPOu4BFFznIK5USEn5UCnCXMIfC
tO9k6MJfIswhrNuTeODTLI1e4y5x/qromp9zpmkIZ/9fZ1AZY4sv+qvIGvwVyM9WCl70f7sJ9uUh
0/et3cUz0YPmXXVdJ8wgmMUmmjtBCIA7DTTPfCQXfGtqa9rUBLah7bHU/iwRQc6d1iz/DqGpJfIP
KzBUjzD7SrZ4lIgi1ax8m7uxj4DMboHWSuhOBp0YUoGhOrCYc0qV4rbitRgUHtUyiVwzKCg9s1MX
2XCrF7STJd2XaLdw4Sj5JoS5luleUuU5Hy2f4LsJBVShZ86HkSgtTCq1e/F0QLMGQt91hq04xSg/
pp3EsYInOtGdjBNmYHw24hUsFm1i++o1+2e7d3b5fhNsqIsm30lm9QVyWY25/ARF2Yan+0YpQnQj
mV8Lyon7xD7NEjZisRuOq+QWByLGpahECohwSws6SN37pUO3nLmMFaFzAsR8n9in+haz5wgAcDzC
1LVs6GD2lSPajc9GAv/v7q4nTdK0kzVm6zbCXUEwMr0/Cz6QZw9Fd75/XYvaYGep0KqqNuLfhild
9JA8ILmv8RS1xTH+47XwDYFfKY+89vr1b+aM4m5G6xjxgRzJjghdej3t+iKFFV8ywNrgk9PDq4Vh
c4U5Pi+4zK1Oj02jyoik37snTa60LoN+1ZnIBxwp2GAyPxczoZw87YWVgqqvJat+1uexnZkP8GaE
Ax/DpQzhwU9FrY6Is8tbndxszr0POAhACxpfR+l/SNBt/nIf9f8Cpt5fIeemHbzMqC/TGUBaPMfl
11HEj8oAuo2I63CjRAV1SRhEcsure9WYFu9zWaJ6NfqLwLNf1eUUWz/VAArgtrvKZ3kWEybFMZsa
X2+sces1At00wo/m+jZUCcu5L23ZKpBNcvML5kFQgoztZqmpJ+Da8mWiLgknOnAHGxoB+k0luaEU
mmzDCIsXoYJOf+0vTwmVcRIz99VPSmEXu7PoLFJ1TzBg1j6Q0pLnfYhULdgQRN7Dl+tHCaMKH0DN
KAu9ConoM3rIAkHXIJXre0l2P4TeX/pT5acqXFEuQ0N06/KCfFwWTJhxMr5YTzeuYLT/uwE+Sput
k6k05ElRdQbCXrv2diDenEdEaahEAEFTiTZtuMo+Ge3SuPkocbnOgbHSAR+GdGYCrk1Zzi7btgNu
uKOq45OdrphHbYmaZaZ6g0ZhOFuxF3hmabs5SUhWXn7HKCyZZZNUuTeDliVNHDgHO4DKghixXLL5
CIElFPbXsDJUB4Pd96R02/CpOtgOYoaivC+kPzqgbISEl1G44aHEQV9TXHs3q77m35/pKohvKQ1j
pG3rC7IgLdB5NfYkV5OvuPc38uYDZiBze1zi2T4oPuISze4OOtZvrtFFKvojFCD4lCBjB9AhfrlV
EdXZh7oC45UDmD2CG/gDNqCht64ZxdShmGZI1umi4M5Tf5z6+G5567BHNzRutms4yqjyfQRVaDP9
kdlw++I512/7DEPv4jM8mr0WaGtMPJKr4MLjARyOCIFVMUc9POguv0hpyLTH6ALDytbv2PfOdJl8
+LasGArxtTZqUNpXyM1JPKasRwGODzmrI1R7JwyikUbkTSXuy2V6iSKtSG8zlSLEfLDt9RIJeKEp
Om/i3zs4i1/1eg5rEg0eOC+wiHng3ycgrjX1bviRRIyxZimPI5IAj8R627yZDwNlmtjfAvKIAE7+
I0n1rLK35F82frx5X697aUVGzbIQtNKaXB+WyJzs5qEpT6G6CUonrCATUHvSbfvQ91N3Mnn0uZj0
hKZXFQtkI/x3Z3JaFlatWtAJT92EMa3mA0Q1Vwsd+uU+z75QeiYBrQIDpZzT7RcHmCiHND18J4/j
XT0Yea4fzsAHRESbtDyfHExRJ9SYGJb0RiNy6Xonxls2VM9tAEFavys6Vw9KmvDv7MOQIxBlWmVE
QlzoOxZirnDGCDjxNkzew9QNXl/vaIZV37ndjqRlYk+02oOu5OMvfGsIM8k6xRYIWI1Cf+yyd3sp
lhitB2VNPfUN6rNIjTInU11VehESyHAVxH8yNzDp7AfgsJefozSup1aEnXIPIkG7uhftz2p0a40X
TM6CMc0i2CTBa62jsR8G4CRs4Kke1XQ90Xbv0x33DtLSnfmHsG5AMdi/aSuumX+NQz0dIcMQMw+g
nC+yGnd0I//BnCAeUNkgOWsNE0o2664Hio7hJ4vSbNb3N6a6Hq5K5caxt1xc4L1auL1ZOArBxHen
M6IJ3j9l4H+WzaOHAKyeIzeUwCO5wtH08SHexpvrHROkIAjg4bKNgio2xbE74KiayFPtfyxnRii7
+FuDEcR+N+41yzRb5ONm4vaLTNrNgyycQjMS0XG0DCZWzKDNwHCgtMq/2nCKH64U5K6Mho3WARyw
WsIijPJ/7Gt0L4s81nV84jCy9Ga1rKPVKx7NO/Pcwhnetrtp26MpCdrN7bryUC9zUaSfPA0cBAtC
pA+x1MLi3+yCkZads6Ft4lV7U9Onc6RNse8Gjvh2hUd5Ecl2gRfu847kupA4X5YAAs/xu66KHe5o
HI5CVVqhR9Vu4sHGh/Wx6Zo5JKwxT69nNTmqEB+zrH23jeL0fApKXbyIWq1EKK/psOQseLwXqnVx
dAM47oCsUzduFNzCASx1ArDjURxteyTId6D3NCauMqCkIOoFwXwyXDYC5xvJ8vYtt644DqM1pQt1
x3csAWEXdRqSGq4iPCO/htj5Eb8r0WCyAGvc7H9/AeGHJA/w3Q1P02kKOvR6aFDijfQI6vC5occ+
CNlfaJwmWEixTZdHI3GtmTCN2OxfvDRL1T87LLcRA2S9oyjG9Tj3vOAZxRHEZH+Vg35MANsFt3kv
HYdBM0mWtQkM3CoTGvD30umODKiLt6/zzisYzi8QYUkk2hxAqeVpJzKmjOVwSYECp2UaRWuHyyFB
D1SY4zDEGboiwSskLK5xVOx/oVw6B2UL8+P3lo7ETx9HOeJIePRUCfE2uch+ELpYaMtKRziL/S/Z
rLO3yGW/1JSu+cVcwZoj4Xn1DTWQdm/6+CuWwxoZf6M3PHRmlHcnvRWMh7fl72oqfQKb0/E7ji9y
yr950IEEh9xLTPr+/b4FSdOtKX+8oRIzlbKtwrZERWn8aWFFBjHZJFrbkS03s7lkXagI7IH1IX7m
KJSkniHitr/nGJtmU6gn4itdBe26bOvmMY/ejfeiBDkmXcPCsV4TrAt0vlg2AsK7QfFWUL1RUJ3q
vNMIq3kCDytv2umq/gizRTy2SdFmwFAxkEuaoUhgyxfjnDYIsFhwSmhcLNBwJ54WMBQBCNbZQYlj
ycjLCnDZqJCa53koyBhFwRXbYL5W5fbmIh59T093cC8/DBWDjOeH109XmKvRgSLeJHM7cEWde3sG
argD/TiG5hcgfoTTZ36qf2r+ppDZtU2BxK6YnXhM44tQ275JR2Y5A1gBpzLOUMUv1onwNZrsc7FR
RUzQtZK9mIJl0/ttFz9sMsJ8I271sf12IbKfTfkQqWcl56sWdtWvi0uonIgYuiEegQE61EHjh/69
+53Csm8eM0534hKhk6iKcuVjNwVOUjJyGkTnMb08LSfX0O46/ZxCLpUxnBVHjaJEjn8EYYNA4jle
6b4Al/11ChG2EH5rDjlP8HbGztekrXW/9OM6nlOWnwHSm9heFivE2RxkQwamiNnnRekigSVXCR9Y
H61YLEdMK4Utah8KvewHR4GvkNZaeNE3kHvCU+0ANM11kOcu37nnMbFv4nzBe5bjE47K1NUeVcrh
V65wt8H77DI9EhruIxaKM2Udlz+J4gHDPWIEk2N1uMngRNsrt4iCxooF6FH6UXz9cykFq+z/EOYU
VVBcDTAsDVaKwk6nFZRAu0oMl4nfi+FbfuAHuTnCncywGPyxk1jWJ5ewzmFvnFCDkpSX1b4P6iuo
uKkM7Q5aRb9fuxxX4DG0PfcoNVi0MsCAP7WRb74aFQBn8+5aZuLzJfRiLR/gwWg6ZN6ZnlQTU1tu
8iSdRoQMbNrBMwX+tuUoOBskl203forelkN2veYjzJSClm8Vn+LwnKF/ejM8LjWU5DqEPrH6oH+f
emKxgNzLiaXpEBTvONfZ+ATd87Kx8fbOjKyaQ7hVVAPul70y2K6FkZLxNcP56+D18FQdTS9LkbpX
nE1ulhUZ91rA6Pc9F7roNLyKr5FqmunXJ794l+c0DW/lqfp7B691B0kad0VU3VH7ZcVYS2DnwiQw
LmvAYmS9g6+3pgwOxUi6wU2F8SlYyzk7m6RrEUrWZAZzoe0IkLfTUgJ7ChU3K6p83Oz2+PXApCFc
Ug9QQRTkTi5zu2JKD4fox7qZcfz2g2sPcA0naNSqVqB4xWV1peM7VFRyEY88wCzahKmb9nOCbXmW
v8pKj8+7+qCEJsqpGI63fgNMHJcno9nTHZLmrhCjEcqRYspXNhYv+IaIvy3KG1XqfzVOswza1i5s
uJKRMKYXuo4rQsNvuvQ8EsFQAKP89g+dEnipiVWAAvrs+IKQkJLJrZHVZOweOWJ2ThpWjETQq0xF
g+Dw2oLfMv9/A89FbTX8ntVraXmm6PY9Bi0CR4lqOQVr3eyvIdlMdjh7BCAZFfehl8U6Jq1/DjTd
cZiSX7Ea56qCsNLFs+fMCz1mNw8xS9sDth4FlcPDzAO6PxwwVL5bCzJDl9cnIw7fTmtXEw/BTLPG
q+C/f3KMctWsUuxhzKkA2r7X5+ETINDUPUlKh1D8WGuCOALk2NPZdSLOT3ZnRV3obEbUJ4swSfTt
u2ySn2TU74886KYncEnCRZQQic5AsfN/N/W8F9vgS2LaRMNzy0e1ifHS0WLZYvPA2q992V2aPiyV
rwQ8oW1IfGjp7aCSB0XcCZmS5gYrHo1Z/0GW1YT14n2wVvR/fktCtWSNWfrA+Nrpuff5ouA0T0FZ
OOTed0nh38CeeVRPP3w4IoHgpRAwjEi941nQYWzK0WlVC+g8tOgVdmZ93S+Sdyc72pp1jUuenu3Q
oO5kBlZmf0cF/wX4ScsAbuRUHG6FcHsVcPg9eKrUKl/Jm8wN67qun94px2fQnhxQwrq2wqeXf7Qr
Hy0fhHq7G13t749oqOQv1BDf2DtsrifUMG96n8/Uy1cDeYuHT8WY6no9xa5kyz0SIf/rcCoPzLjo
tHATT+tSiDQu7SQFfkZX1IPtpC/gQri5LlNvVRevo8074slPbYSOqZ8rVb+FbGd40B1BfIdc4DA9
fl8px95bBq5vjW2+YrgFn7Rfh7KM7s6SfuKUxw1WhHU3+uKcnscN+qAVGLFf2YtlLxQftdeLG1fx
U62LtISNFojKP/RZxj3r0SFRWY8celk2AVP/hKGWOTsDzXnL7Z0qv/S/Zjqj06csm0dRtZHmDiF4
bdUfP+d0qqlks9MhCpz6Wj5Q0Wmwau1Y65hQB9xKDORPC4pCtRh3aZkCEYn1oOwhaHfh9LMRnMY7
0gc1CmbkYGi8Zd+hgtMyfXSTZEIlH8rXuXOhzgXbrOXbcFkUvbXqnzhe71LIUZ7eNcyQ4YHPKy3T
dreiZVSbvGx21KKzKDh1Nw2Lsd+kcL0gC8lnNzVINQnDKoY6MIjaM7GiFGbfvbl09z0kLsExpVdr
Q4sjVxQ0pbpX7uDMcDN7SE3aSwgLs07aaf9Ms0b+Ri/Hs987eKFgYQsl8bK9mTc1exWiZ0MA+RfT
hZ+KEn84y6A25LeZ0u/KS24GYi6/mOh8wvpZlYeOnEHg1SJF3+n+kCX1htS2gkJJ8yI1hVdZLV1M
M+NC5CSapzLcIgKNB1Yp+UVF7Y0apuCXgduReM7mEbekWB2+z2ajaLlJPM3Q0f8GFUOK1NJrnkQy
YHOu64Fn85RIbh/bReg/7PywaStyqhex+LCqhIJtRQIHVi8vuH7+4CghRlh5sMHUyCJE6Iy5a9jb
V8/FsNEdpvUDafTL1E57f8g6EDoz+9d73qheVGyKgEE9fGf/4pEF1d1nsJgcWZQwCppx6BaaY2Td
O8lGdZSHh+b8aezupsgJFerkckUynb4zm52YBMMvIpdzGlBO6RNYQoGeE8REm/ls3tRyKWWWzIw3
IcqazjQmTgM1XgjH71IeUFpy3H+1yuAoWLujVmK8iZc1ca287NId9CRTElS4p7p97H2mQk8kF/nn
Aa7n2A6qQghNk5GvbLSzJwJ8RAHgmP/vz0Kapr/LOCNkATecXSo0E+Kmw1dV98VeX0Ai+dxPVRQE
f+L6ebA38FPLmU/B3qkUwFymcpvjPX1ZpncF+UQnw9IjMNHMxkutg0i0F7H1fTornShJCNvOgioY
DA6sniYY0zdhHUKpaU20os9AK4GHzm2EcV4zgTRzs0nJJZ0fJH22tqlCtzmla/NFqTfAtHQTZFIv
cHIXcuEtbAVOa+BDhgeJP/aqb2QvTJig+bJY9ebTxP7ekFlnzIkBc9gusacvVh6KF3JpOsWBzYef
8Pkzcw5E4xSEjlvY6wHUI+XvAWWohesOV5W+AMUJBJiINTCK7hPT/O2Z0TZyFWyMTe9ykUlpOlRG
vxTcW48L08KUZrKD+oRVl5IaIZz/abT7rV7MRTOCD9RGjSxW/RhR6LSfKgg/0tb6SCVC8HnPnP83
L6xn+WyoL5bs7W0ZzX1Za2qFwGQHjuFpiKCou7XCo1EXBhlTlbuPr9omG861cZurvHU+LTEG0Pjr
tZU4iHCaZK8lsXbsJZkfdsxni99cAU+s1dmyqKbbwaaFvGXPNiaUtohddHeka+ZrbnRp8ZSvfyx4
p3+rYvthIUiY+OX6Leb/dWfhLrv8lv526x5r2dRaP/03P9aG0wwn4TUc314Rwigm8y5VFygSuBk9
gFD2j8ytqyqtiV1sMP9cEyOfABRxCHHtKjkoTxtzLeRq4GcznFNP7KilvSnjC+0ctDpN1qJEaZBC
+fzClBYByj+Z9nbqwe4eSvY6k6XcmwNdMU7bduMwNsCr67f3tIR8oGVm5KJExNszdlP0tJxR15WU
7pGvbHCQ2hqfzU8e5s2MfGM2S6gwzu2uc+Igy/UaQzUZttw+97H1vNuy1Ksl2rj+ZLcISntTEBpg
bekJEomK7axepJ+nJwEa+JeKCLAMl7O1G9BcHYTnJ+Mn06h8ObGPUTT4I9fzw8XylxsmU+9U3awB
Kb5IIiCB+LcphZI9uRySHuXlV/Pvx6AdoBFqfCy8Ec1SmcDK22NfLUWKuxjBkDVHs2OmSiDrtp2M
WKaAsfjImJsaiopc3kFhVK/hgb4QOWfjb60VRo6xDEv989I1MTZJ9quBQ+N8Xpff0UpcVUYvmndd
7E4yFzQuMqC1uJMqkN+mpMseXwevN7bpy816zQXO7uki0VugSJH30WpSmJo6vDYM7UXTK17+Henb
eCa/lZQ4T9TkZXepqfzCZwWUO5SO9MVH5YOICUHGN4lJIBIkUTvUXOjzqtaApjFXeXhZLwhErvrw
VJNxIWuwBcEuK8VOshVVUDDt1clhSqm0XumaSNd96T5ZblwkMc4Bo53OpbBNxFjQw7pmX22hpVfk
iwM+qoutynzskJ+lqIli7EfLgNr5sqBman4uF05CWYHk3xPRURS7/iIr46o9AQsTClrZJIMvqajO
mMu+vnDK1s82PmYTL+oaYuER4tQ/R31Gx8bSrPsXMqD9aRJ9okKInOCOYIKAIhnK8NJ73deo+Zh5
SM1egWD3Cwl06h/VlOqPZeF+7J+jg1YKVhwSBJE4zbLNKPNNRcydtylbcsnQn4l1fWovImKUOkfl
SIwVKl16lsT9HmxV3ps1WE+AsJCesOFKH4yxVCq8FuBQzQJDFsUUUdceJu33loQtMCCbrYwZt4CB
SKSEEO55h1+bTit+qDc5OzN9aUk6xvzo29tkcnULNcYjHm1tIUYURu859zFluXmwPjlQvBJ4xscw
ejL56cud5vAb3H03PxZN+91jNBT0drhmy30Jch19R+4CBq5a30CsZ/F6fXTCGgMfktR2fuCsjHUZ
97PP6HTRP5R1tZEfZf9n2VNhoXdB2lw4S6NgfWcpkqd4lluR7QszL8ve8Zdd9gDZlhfR5Iz/NpgP
qh0Otpw/Bj4w0pSvTFqLDw3nhrqHSVo58RL+6MA1lF9ZBDwpraYNglrU0cYT/UwmZyCjwxnkcy2C
Pr+xjFVCJ0Tt83xz+QTrPYBbtwsufgfHzutmsTRreuEDfyfBjwU4JyOaHJsIez4EyV/M1QJsV622
+p5NRB6VAyOcalnWAzup5YMhXs34YUGxwMZXXih1MtkzpavZRcIfnTa0vs2wcsI2TlfxufFZXFg7
uopG3HNdHjbhCYNJm379MnAYMYuhqaYaPNCTPorzNboPf9sIZa1vxHEadivyzXOxHLwq2zp7Ovqu
OWdsaLJbj2r0t4BhXIkYE7Re1/HChnlLgeI494za9QYwjCCOke3PO96kSnNHgzCK9AOdwkTXyxb1
UIJ5eA9yGoZ/I8AT630TYk0JbCaU2shhiucCFXVPbX4XznhjIjrvG6mMxaDIdNlOvNwkL0Eond7t
V0HcX3pvTs6ynV0kiEbVTgLkRaetTuiIS2PckoIONbiZGmAgIy5imG4bp3xGII+OsZDgNrTcRvvK
URvq2Nuz7yGG573mmplBsNnfpX9ARnPl7tvPaKN9Y6EbtueizNB2CubvwPt1rNXQKwFgsCW6A6B+
awNoNLPMNHbAAt3gKg5FU5fRff84N69ZK0Fd7OOc9O9jTROQGr4rMDdjWo+FTEyuZ0Gf7o3Rt2Pu
lR1xUuxVRiQPR/0T/g9cv/lgtsFuKesToivBlzbRNhkHVm4m9whBdg+yGaSu71b5I2U3cYQZOSXx
H8eFrNrFaBvlUd7JRXU8Eq4e8DDPH68XaeYDuTKe2oJpvew+E4yLS6vlIZAl6c7n7f+WoqWqBsRC
Qre5c7CYCnKzl6f5vxOr8sRDzx8w1SG2pe3iABlbdKcsAFBzqau12o6TZxRH2soTNScz4oO9QP+3
Wk8fsqlBe598hT3YY/HMoKVykAhI1uJLfevv6K1yaeHe5ZjfTIAvCEGbxmMvHvE3KymvTtA88h4S
vjrwfScKxXuJlHomh00nzkUYhMGpt5+9LF2sWEouOVY2sWAMUsDSyNxpst22r9djZfEJbfCdNUNU
GiLzWzKrNhS1jN5pMM8WKj1LkkDJULzJBDlhrakcr10Zw9DYXBiwqitP1t1izN8MQ8+XaSuVQDoq
5VkL9o9mPGpKcaFQVmKkGRiWgtWHcn+irYyle9d0cRufm6gIs1UnxUYSFiFEo4y7RY1/q6SbrqrE
7PwetQ9JDs4pnjIjriIaXSJrZxf6VmUmFlvSlg0JKtFcZ+a4krEd7HZzi8y5lfk/m1bFo/zw5Rhj
hJPBmszPgU/i9iSQjORst7b1SsqXC0+VJ0U5ug9XZEOiteBFX1eewPqqZrIgm5BsbJUX9rtr4xin
OESJ1z6xVT1uAmobiMJUX3dW6IXnx419NSPgEWIWKMq16oHsjoO7ZKo4Vf+UYKEpXYEWAVYYA8ot
v6K0y+JhRR66TXDXeRTaWoIqtmzOtOEf7qSH/Pq0jTaUlrIbu5Y5lz87ImZxK2UFatuYRmZpNfDn
PfRD9EBPSYh01A6+e9PBhlScYweUMG0Stms/L09cnK9vQOmx8m1776qrJcLL87rF9TtrGBuEU/rx
SRCZ1cH0DdLI8hVVlQCBKauOYMcib9vnJcV5SB0pnhGYr99+TrKcfNb/WHiDqH9m7+/Ci2Rt5yia
uRQl644KZHx27jhpKmsIQKY/80PlZbZc8xtRlLnh76f3eW8wsgWBdZx1xPHt6u/3/G9gEAyrzjpS
C5tl++t8gG931gk64DoybnUOCIdH1d7rtzHId7s1/pfx5PB8THvQIKWuuZ5wWiHiPxejXPQE9enn
/zI+jzZkUWqZ7ModH7OB0+vlQPiwjEFaBVYpfcuWUeLv72a3g4xklRMjNHS1m+p7BlAmEjzWQtt4
XTCupey1sYeUIiRjaFQ+ESImVHIopwhHEZeOcwCa/thpD9YRs0qnARqlORZ7Z/8LNlmASfH32rRG
FNXfC9Uh4rSCsroga3YTdYkLkTYDOqKSU2FcjeAA11BW6Z+zhQ1naNiXVYsLYAPcxzvIJYSzVSS4
j/s9NqMF28YwlMi+O5I7l4CeuypdAOKxJ7tcIiX9Lm6dXlxn/HShfrFFWyyUZ3QgCO8Qdkpz6iIX
JV4CYt1bhGT/dx1WvO2+BFehnaAsnjrpRr9Z/Nd/GjW07nadYFddGgS7izC05PUw0ShieKz9Y336
TQtAp4dOSzeHyizIY9X3aCv3HthwfVdE0MR+bQbMoREsFMabujXL5jKjeq9G2ZMebKGGlrVhyozM
7v+egMDjFr9MgzwyM9SBf+EQRIhDs6aTsEgFhJmiJzh+tCWOulHOUfadKhmgKIpYWqV/5nXKTdcd
Bw+MtFRYdjDujOkVA/aQpoKbfpOcCdVxTN/PVkQT6P2psthSNoyh6dA3JQxNOX8/RAa5zhaT3nmC
0GNELFPBpjWHWycT8rJF97YgkgVVeUd4m9plJiNsz15oOZUuMjnSa5n2xKSIRvqUiJcteYSSRHrw
SKpvO98ubzzfpTE1uUTpBTyGNoAMAuDXi+MT+KlgNjecQSnL8H2/3V/bR1l8FccbsmdNIwg5KWZc
AGkHPyh3jpBZ0pGUEsvMUKIGQUU81dB8wYWX+q7imNpAWhOMzBNJLzYCGKQvWiVONDCVKBSxAB8r
tIv11IGZqcvcvE3LtkYDIMBoO0MkLCWD/GuVu9nZFDGjlFOsEaJ9frCbPtKHhWI+EN7lus2afhzY
/Ygu6IFKyq03zuyCFcOI7gNgtDVCvjtNWn741XMe53curLA5hXi4TaeLhy9xJbjSkCeLU0fKaJ4b
GQjyrPPaqoMNHoDKQOL/Us5rvCLQa2svl+zYGUhQj1q+GShNZke2Mw5wgBoz/jmq6Qo822ButWH2
D6IrQ97wowo24qF3Rk35Y9ffuCrVtAM+5HRflioX+INh5sQA3FE/ZWF8393bL3/slnB7D75+M+Jv
7DGw7cZMoo291yqbvEAIu2vgoKBYp5TxcVzlk0k8siSjd2/SUM0kTYSmh4Jwl187hIEHUW3UZIYm
UPNLogAOhuO/0i3o7TYT7/1qLYoSHEcJ20PRpEZCyzo2RdxFLWsEEeec3UT2IebXEw3aUH9PuUzH
Nfz4a1EJBOeATmbzn2l/67aoKobCaJoordb9PtBDXRsHeTbRCO+6ajSquVbzwHjebf5ClM9GiXUX
o/pmFfPvWR/6yZRedU9I7u4aAYS76uYvQQmOvO5gBHtuDg3hh+704mgIbUVHltGZ2giCByTLQsLI
AmFbR3n/0lB4F8ECn+HPqYEn9hNcCG/k/7JZVqIsk6H2Q0fMQf0cpTHBxLrN4WMw3ZQV+4cB+QQT
TxdN7v1zeOtH7UgDrcaXh4/C5rehvPg1Wh2XQJN4CluaRW4L4T6d6QaSojFNKvZ0QLNRKiP9O7q2
vXtllITZLUfGgxeqILC1nDapKwQxduuApvi7v+E1EspyamCnNCZICSCeT1NZ4MrbFvti9tzUMVP4
meApom2Msa40UrlcJcr0MZ1Wnnaxs4waKDR2fba2cBGNRCCmcTGX6TtxsPf6wMiQ/G72GjHR2CP4
qZaYzKvFUKFdsgb4YVU2D78xDd6fvfGPV3l1sb76/uxPTxPB4kWMbrv4X1HZPmTroTmihpS4gn1z
xYxABHU8h03qA35qZj8wwn/0QfbI8lLHj5kpcYpmIiGW/WqFQiJLQZnE4r0gS+0APIhGk5qmB1mR
6SYfo2B94JwK/VcLlvqihDJQSMvCCm6ppK27JDLFJHAaB2/9UiVbg9IbL+B42zLAvHUvwwoVT3y/
nW8bqLmyaqzrDQ75EYnwxbQp3xUhfhpfdLbM4m343UkpuzzvypKEus1dM0hWJd7Zt/R5SEMMymBw
S8sXSJ4der0X3hDRjvFj4itsqWPxwZrgvTDl7oo8swZey7JbLC13jycsm93RMu9o/z+snIDQAeY+
7Juumqz/e6aW+KC8lhoqcakzxXyDbNR5BuhzZkzDGGkyRgUG1PmTa7Rl82gt0NR8Oo6F+CLHqzsB
/86DDUXFQwu2kkEPUr/3s0NcP/pPIv1aEszUGvuIJm9+KJgduLKlszIAJPxKwDk6TY5nLboGUB3J
DAD8H/he15rAXY8Ah9P5tZ60UV9y5Tj5ORzo6+Ib72oALrtfzb5fmFL7tHfti79akcfPKU+Us8j0
jrOZXs0fAipoZ+tq36/Hk1zcnADRpDS7px7tX60HBAJ+V0wi1+RA4LdaeWoTy21X/47EuK4wDP30
w+2K3XzwrC77Lhvt5m+kqbdmV3W+nr2e8cID8NDyIQg7H0LUKgsYJhoBdodCkUYz50DaDezW44W2
WD9asvbwb1h1ZPmobHBlKo26eya6I8utQUmqQgHGxEpqFGIsFtIV6gXrC5D2ED1ggQsabygDKQgE
99iKgBfZbu8Rv9i3yf55/tXbr/CPGDkwkalNdUaUej+9IPBLfv/2VptPNiZ/9hghZyaxk1hNcL+J
KUOOAjD7gtiBpdEcSFS8/TeY1uzQDkIuHW/YuCOj+GPmwS/k6SBvzn+Xj/n0fzORmOdsO76XQxyK
xrWO6UH6fbcmdgKEfIGtrQI2sXQMeKDbXT+EA9fwDQFlfHiM4c+/TAQoIrDp4qPl3Ht6bF4pVQiM
VVEtjPnnaHWF1Hdbg8Y0bQlMQIswNu2bCkm+Rk+n8SddUqwZv4mugTH0UiTd1wdTT89A9KwKt8m4
4rXtkqkOn5M2ls9BS/e/7L0GHlx3NSaV4zkTG8BMlHN9dRWg0/UTUtenkCfKZyfAQ+B8Firf/W+g
WeqlKCkXnILC4ydfBtsaMwuQDLwN991rY0HFdmj/hc9zpRmzoa/szJoFJ0ejesozuVLp/u5RSLHY
Z7xuyjDdvsUf7J1a56g8IUayoWVUI31hVVaIDyhMOLrymsL6eU+NqqybRHiJOXD7Uye36wp3fFNR
1yUBxfiWe08UInJNrF5GG8C9BNJNfRFkaIDBbI5lXR5afGpsNXQ5RUUX4WQ4P0xxUk0wG3Mp9wYB
rxag0jaeb3ww93VcjHscSp2tSOdgcO+dzf0LyFVNDtiUXRuwLTn51fAfas72/GjOWTc3tLIpC5LB
oNHDDlmczSi3dDLLLc95SvSwqWXe04jGuWc+gDfim9cCdjePPv+XuO9jlw/YrE2PrJTtRpi0ZD2a
c++WWwwRZwYhO7aN/yS15ZqvK6F7Os7BHHgBxcbL+ocAhi0UYeF0UZ/Fe9JAEGK11dBD37FEinc3
DNnVh2fqA4Z2EMdHZzTi641VI+vmPngDPizhvPXtlmvhA8DunTaQZrWA0Wb79azWDpQF9gxKux4f
A0jFrVi7/q/addw3AWDsj1yvlBa/qpVtCzJifnImZbO6eTYhPTY6deTNJSZaF/ISGYF5jr2cxqzX
vlXyHb3YiWH6clhdm5dzWZ+ixtlbXB6+qOQUiboRqrxGVZ2mTiWV+7gugOwf7ZdQf4QcXscFZzZC
eFlLZB2GwfYEhMNYG67VQwfQo9aaF/T08TtSwpz9prJRzwY3CvaFnYUatInrxUf2z0vqYCXJqEyX
Dl7hVwzmSfwppHSVk7tJiI5Y/4wnhPf46Oh5aqlMQHkuj5TsQm7ZtWgA6kG5/XuSx5lC9lj7ohEl
OOfUUhMX1j9IjEJX2ppchoOuPfHWJrTHyoYmiAd7qDGf/XJnLWOY26TJtEz26zEZl2jXRAebWh7K
q2SYPWdrmsVyxnSLMZJlXJHOZEyYRjhECPD4yA1SAJJASMDzkVwnXqzZm6WyYGxbw8xOVfVUO+oE
+UzW8BkaDDI2suV6NxPvhE9gC8IZmytUEt5LAV8b3wJ2Ml9HxLKs10FK1eO2ozNMcPWswzDtqYAL
nZ4tsXmT9g8DDyVyM9EoZXu7L8jW4MdEBgVy9QRljkelGePTUOphtyBWV/JN0MdFS3vqWyaGvaTi
7MaOBQFHGw7p1VNxgwxjjzEHPdERQF4MiC3B3O43eyaE5Z9rSDuZNTMv5yjFqah7MLcWoV6xwcmu
gygXNshNNe48MntCTmL3mmeTEztax1gFGJcUgA1TzA0GTJGmiz1nFkikJY8VBJLuraCD6AhRJBeH
gOjrbRZhbdWujZsHKhzy66uqzTmu9wn3qQcLQ2Rzl7LTKHMguGbwjrGr06pbFcvNNUwC8KccWdKB
MKlK3BDrF+6axEEsx3nKMpVPqR6onHu+DnB6jffKay1/wZoP/PuxlCh7cCEDuc7Plng3Bqbz94+D
09s6UNmYio/02hWEJ169LOaTSSJ9f2zqosu8XM352Hf+yoT7nvg/dHvI6M5r3yW2QVUs6QnSf+pb
U25mqZ9FR35E/jtBGWF1fwvZiA1mxrh79VX/pw2zxm5X/86odWDeHIOZjWvRP6ZHMnP2+6plBrKe
t9IyIPvYbthlTUas7UABwoHXOAeYPK3V+eIKAHrTrfQixk0U2xNyXHyG7UI5jYjfOTlFybpx+TyS
mpDggFzPpedFXVL9SGU3nPzUBu9oje2G2Inf2YAAfONycJGTE6bkoQdT/cIO4n6Hl/pV4uWzTByr
GmTq5+p3cVJKbpJXFGJ5TaYlA5NB+n2th0NcCLHf8YDL2WcUv/sowxkiDYtC+WDzhlkNouQFaZOV
wlin2un2eAjgM35yrxlVQDMQm1QB+dvlb+24F+cWyn7OY3md06gk636+GTxEONIr3CYMawFEiuBe
Xt18Dd0U5tYswuhb4rRYu4q8++oKu8/2k6sTfBwfeR2ado+yXjdbImDYfnXSpX4hR6c+aQUnOgLi
+TZbmL9lLrYnr/CENlIU5cCSNBem4Xcma0dQUNDeiyC8yO9yDKQ5qAZxQzipTZ8VXfzr+7Gn01fK
o7UQdL0htc5LC+yq8xmQQUJipRn+jnCQ500PT4RYeA8dzLxWqXLVoWKusBqvBodpdyDs2tMatKh7
59U747Q42g8SEya1cmtNPLQcWrlr1smHLrSmi2sUcLJPW51nGqSPyGkyZ+F0mJuCR0/wGfv5EDhc
yEzEgoozENV2ZxuPLFJ3GCBxGj55V6NwY4tu/UnjkBP2FJ9Ngo8C1odxo+/FuK4w3wdghdnWXHVh
c8CqOQYW8Fh0nNbk5vz4eJocjicMIut3B6LcBWmcHISk3lFBaYrVOYpNUjyMeu3x8IVyeMwYIfFi
VG+0HEFmCcCKjZcxSjLI0xvdG9R0NuzTA1FamUCNGsqnte7KytsFEbN1w6nJoH/pKoZA44EqY0Tl
gW+I3Yp/fZGrqVohcb9BBE5X56GVlL3aqzgR/8Ffom7CgDXjisW9gUDVgVAICllyisVT2xXleCiE
qcCco3p+2woJRYrVe1hcsBKpxDHzMdy1LkpqZNUpejlG9rsQH6rxquyHxOdcq5C6je/HaCCfLJkJ
4XW3uxYbu/iNBLl7FNMiROQVY8FIm+zr242FZlfeNtTdg/nNpVT41xPVg8dy8E5DgjFFSF9ozJ2R
ci1VFXGGfk7yxM3NlDBZJOssucWdMHl9uyufYGr6DbCvpziMx8Yjska7dgpaS8BchcZuJWpx9MXm
DeWPeyepOQ/q0sJ/m4FYf2UUF5mC5beD5jC5KEnGZqtMUMhcreEwIg2pFabjLEXED3YZFDqbQGQl
2OllUsOM+FUGTDq6ultXVtz05aWbe/kfEt9u491/Hv0aDYZYCPM56xhyLJqCPpwlx4AydlnLsbiC
4kgOy3CC58LmPOapLz/feZvVIffYCs1oSzcKrkrlZrcq+01Je6a/r4nDqlVBzuFC3nKqSPzNxS3B
vEYbR1Xu+o3fwffrR2HuJl9Rrzthlege5sEIdYBaHY1RIiX42n9jVi2p17gBjUU11WXbC0yeP9Ew
YmeWtZ0xM3ddP/TC3BY5I+czJKjaVXjYTB0icKraWMnl88Ff+/t87tt5+aMfVKy38rKLtpQZNVi7
phRnSgt+JhI2y7V2JPq2HM4kL9fEL2Iyz4r6xmUSQSQ20VXFyQULQmhtq56CE7sYsgznRapBQ3tb
m0nQBO6GwRnbM/Bc1IheYCI0dSBqd7fo7vxmL03q1IX8mthpHrgmkgNoHuONROEjlE32WDYvgKN7
1RumLYSDXSsPlJUAecD1KryUPK3xghkvtueS3zKv5mxhjD3NhgFWwUI5usJvcdlMvWjrJFyzQNCv
MN/Dlo3cn3MfZKKQun5umSD++9BVPQvt8tZ4qU8MjN5OaN/XoQiZAdtBxs0G1sRJu+5X1F5FrQjj
SIem3YUO6D8W11PTmka8ZiXvkjFDdwQVcQGeY+WPGQktxaAlba6NGdqcs0GQ+ZFXKRJjP12r0CKG
QnEaQTnCVzf81Rm4FR/U9CFIrBw8hHgXL54wOmPuvROTb+9sP23DLLC+/iN2iip6qI5SGIZ33yn1
5nbaTQvGdi41Ye62OqBof+qRAjBA/Aytb1zvFdLtBVp9YETh00zDLUX/AR2eHSnVeIsl0Vr4Qylj
fXAffTyk4x+hCkRLPCGEqDeMEE3HWzY6BVOwRBzDj4VnW2CmLtIZclxNcEVoT6g9kIYaUJMAyXTW
HvubSsGRW9H8bJV4jiBMFP7sRZnnng+nw1jFuM3rh4F6LBxkia+8LPKn2ocIzmmd2WcUe89u46T7
V74k89s6Ag6DTK0dYdBt6+jQxUzwtEtuMTwf/Xj+3MU4k+siGtUWTRcyJ/08t7jai6+M+Ma6br0U
BrIQ/d61a+i/o9VvOPnaSofpdHdcEysi8C7uWJa57uHamJarvpPVaffbePca9DVew0tB7d37LEUZ
h8E6+Ua9/GhkuCc1XzD7sJQ0PoB1yVCQGvvdlhNMK8NfvojKQAJoo8ZGjDjzKzP8boT//iENKoP0
Ysj6U8+V+3AJRnUeygJE/6d1kOzMGEDSzL16trG1hS2hkWGb4IBUMFSvjTH2M7msiQoMvFLskR34
RjXkcDcA3GyreY+7/VM3gHTzU3TZKIpKKQxyUccejQ7pSBlvkXPyQZSDYOs8yWgT6AIBbT+CVW1J
sWHheiYJRU3yxrD+WZBk46vuaIAF/4scbRZpQWdHkZGy6kXA7uVUhXvkDt5l9bRkR2g6NkQU3vgU
HodyMXLJ9zf2SocS93D3X2/kdPdI5u1oanxdA/hLDYrI3sfnpGAJrUBAba9RJUDBiPDEtfTXpYy2
2Y9mh138/0pBt4yZKyi1oSMQ8KpXWWDS6I2HYof03DYf3kUVNNCujOYCiib9pKjaS3og4Qa7mJy1
S/0wyiKqoyD4YXg7Ika9xDUkW2gyygGGrxEBT4r9R/W/Qx1JZwBsGz+AVUKcL8GbIkgAdyAf5LBa
DhbyCMz/vBCY4EWbcluJ0D9aNQ18KJnkq1ZJKJelRSb0VF/QF+3xkb5Zp27uQI1R0a7yTlyUPoh0
EE+wqhpLT7dgQifUK/tHYTIg9DA8+Oq5eppuLQdr2ZmxU1lnlUeeXOyG0QXM6B+Kj1XIe3Iutcel
BHEcPrSQvpD2SnBitUveKgJGRFCknxsJ8/C3URqrPNooMRE+5QZ0XQhFqV4ITXWSzm8A05UM+zBs
Arfxi9aOZBjZMC1zKhTjXDEDuVrNMe9EpvMcJe//AyfmNpCx0NQcOWHwbjn0pdnJs4hh1ZXJzo+W
dfGFFjBN60U1SwsW+LVNAd4rSXwNw783b3h784Kbn5Oem5RyYmXyytQ4l17MyyjPpCf5afnkAAtM
DfVC+wv8IVA+p6JP0Y3euilQfbFQYmtrDusnFpIx1uz1DVHj0l/apffO4JXheNzrw2q5VTHSYlxb
UuSTLufgLoqPZ+2J7RvRcLHRUeCZrsy6Sujyq6WuCLV38uqRSTa4/PiCMMwbKkg//goz1yxtM3ks
St7GU8iPBQMci14d5A5iRVqDEok1JllWtIqKUA+uLnJI9jBZ2+39NVze+obhQ1rAK7zp0ngt7pOX
or/TZMb/Bqli2tBTJHtfn15XwVVdbXkqLxLxGSNJtwSrzKJvNG7uS3v1X2Z7OsqgoQhzkpDEH55D
gGXHgfJK4adIQ5bj9JjFYylwfJODfM7PEP47+wMmUKMlXee6roktNRVaSHOJKGALkFNMc+KIJBa6
u2RWnw2Uj1WZR6io0eVb79YDlCjabEanEWF30M213H24788kf6L8rqPSMMD6D7j2TREcmRjYc9mL
yIFLMMWBtAQPA2TIZe+y/wql53NUvIbupUZ3bm00sMsOKZYw+jfvQRdN1nv9b4mM+mV+C4LZJkmT
ltXqH16GYUISNIqe+iMTzlrzIa6TbFuJ3YNGUrZW5QJn+zE+C5bwBVmZztiHY6Vb8WzoRaPnPK8i
0OQM9LRVIFHbIi9+AJsxtxMw8z6/mX8szF2khwPz16TFkphlTPmKT2VG/g/tuZfkq4UEb3kaIN5Y
piENl19Yry1JTr2bqc3RpUvPZdlaCApnNF1Dj/Y/cf3M2VUmNFUxUgefQDpHrP5t34BVlSaZQN1N
DZxXO+51jL/RGep6oC2amexHQKWsJuj7tBF1+gaP79ANSLjKQCi52IS6Tbi3yf+IkByqUW4nTFaM
FHBP79NtyAIIOUioq3wySh9L6QlhUA4wCgv8F/Z6b0kypagmHTpUxjaUJ2ObNTslPsPCmkBJ0XG4
j6LfkvgVNI2CwVJDTLpROOiJ2omwjlTEahxSehanX+JWQcH1QQHx9q9aqdpoumNIYlukr7En/abN
kCWdDGO7mpt2jRbNQIg7gD/WfnRr3fkoAcsygkDQLgYTgexb18K29eBG9g7OkHumKI+d3ikYFB5O
UjuJbENRg6ggoZE6Oh7XsAcf6wFrikf28FNig1tjOXenLyVLcpymna2h8WeqfkgABe8xowPCtfSh
kcXcOto+z596EIZjiivbDe488Bfo1wKz+wBoKSk5ZeCETlwf0fNNZOVoiSDVEU0XZ9HN/Fm1zpJC
nHwvUWDDsjnwN+fqhHhtiR5XCRZCyzbpUM5w6FREL/60vcIAKA47ElLioim/34fo3w/Hyz2J1Nmz
9iRKjBWahZoWtmHfHSvAfs8760+eS/IpUb9nH2sH8ilTMLzxgEtzmmjRVNpqc0LsJs0anF3i5Vn9
2YMoKZwv712wP4TDNXCrzh4oiklsxS9RptVct79433TNLuZ2/d6g9Vxrm7dkwhrweI+jPmEwVVJo
zO+JfnKRmxL0J/W6FhoAoAAr/WDuzDit9ik3yC9RmTZ4QP+zAsn9CZtkbH+1YAa1FXp4OSgNBgpP
dNgo2Es0uMy1AA9eqB1BZAfAJd1pRXvhPRvhzOSQGZLO7QMmB0NQOaipl6chwnZqCturUT8/vy8s
xZgYjPaM1Tx9iABfD06RLHySDKWC9KA2BnwuX64OgTrENAk3eSlTD9+tH5P2Z2krNGWSxyl14diD
jF/TMMms9Qc1IFyU1za5T+/Iacp08RPeGWIC5FOymTaIvYfXMwcwmVr6pt5WvakBqskRtDH1ceaS
hF4UyVxzTBQ1adZH3fPhq4VGuFvhsCgo4avrsdLOuG3Apa2tyEulJBEeOjl/4sQa+KOibHPC6k+e
XcML5keJurEOH1FsNrxQzKwYibdst78Si35vrpTycsZ1YeSa35ex5FpKLuvHL0e5y10j4+P3vLYE
i+EWUkrMzZu/L0C1Hd2oi0DQL7NV6r7pzJ23ymweC6Zoim4C8mcD7ArRgQw92TpnmprQRkyK8v4v
JzdiiJu46R+BHTUjnpzM4HHHBdJp2GmOV/mxUPmmBV4OFbhn1kn8ydIBKzKK+lxEDHcTLexxIf5V
mcGdk1ZP9z7iy4OiDbDGr7/10J+e/ZUFmiD7BNJIMRzdyz02t9hSFWNqVXgiETwFCibNh0DhBFwA
DHehdXIzdrw4k1XVE39+fulzcKkMrRqhlNtcFnh2+GFnT5M7NaASRzanP2LHNLT575s9kn6tI+MG
9ciP+JIJJYq/pcKFPeX46C1eOTm3id2izNi+ssTJU/bSV//GM7Y+GfgpRH8hHhmEG0lRn2jwUtl1
MGSKOVqZaV77o7LmwRnsvPpgjcNw7gFc23t/qlgqiUwr0SvHaF1f3pZ5OouTgaUhS8zJ8tuVp2EZ
V6MikuXVib7Z04wOFKzoEESZtPblrYHKenI0pP9nXbFxyvHRCgqYBO6bQrLLP7pmBUqPk+CF+kVS
dFVsmWUYh8kS9scLqtsuRYpxod4wRhDYttMLr93VsFNxooY7q+bFCOZaC17tQtkSJ/TcZp8LLb9R
iFo1lpM4PbMCo3dYGFRuFV+JIiKC8f0U9bAn9hGkYptfAFHXaz0CfbvnJh+5iPX+icHnhuI05QHm
wKvy/inUywviU2MIz5NMZWkjYqOYeg9YTNau32jVuleL/V9lzjslF6BeKjqT8BFJUZ+OBB1+jPRU
NSZ5plIljaysH3UQllh+Rom6ftZ4GZbb8iL1lt2ULxU33j/ltRW5n4pqxk3t6Jm82VOh3SRuo1NE
n3PCQE39lCNXatxxWQgpkhewndfWOQzGZeQdmaElF1TnBGGfT6K6MSLN8KCwFe5GcuNnh+n+K3jL
VoNWPfJHjwPX6BvURUoD6Kzkexj3PFA6CJ0+wUtVZGrDzW2XEMK6zfvwP5JIj+3cepkzJzhjHNdU
7/NCj/VC5UnnLgc9eAGXoSKsUrnActaGnnTRHP2HE6Zg5FPreaeQ2itscBvkDCqr2SA0wDyFA4S1
JKlvFaG1Z9q6HEg7CTkfYrssGHqam53pp+iEs5RWg8hLRjUuV5Btr6XND2fne02FPSE8cJeoZdP3
jaEbknj3GjBDguABiQZLDBR6vw70cSGaNHT7FG6wiq0iSoI1XJji5TXBMIrDyaPrDv75eOYNoHyQ
73PqJM/4AGyzBTpCi2JfqBOYT3NFghUEjCvqK2eyhJ5D3+tfPro3q9tfANArbi7QFNiPqwxUAT5C
WyN9ZDs9lQ82omqWRxWztb62Uxx+WSekjBbqN+VcLb5pXnv73VcLJtexR+eap/GvzKPBB7e/Jvwi
JGBc08D2eR1dK9J86ZpZFUV7iRZuGJJX9xTB3SCfda0oQa0lJbRhYwsWV5D0X2cKiI3Ht5yZOB3C
uCKMMFpV5NShwmn/MIC4fvXKlXEAeWukRSntIl1W7Ui6Hg6GEeEjWd7hpSrkXSWNn1qQPOSLr1Dv
ui3FmepFJbD7ONRd6dvGDmzG0RF3gRUg5VFN3bOsz4LQTj6oAs5j5U+TTjrXOP7MreZ5ILKKhkPb
+iCf1euzmXo9nFARBngnUvwBbE+u1pWKLXWcW3CAt0oZQ+8YrXNXfZXaFFmVZt3EDoTWArSRWGpo
cQm/7NC2Uu3tB6/6olEZiIYd2xbF+ri4q7d06WyUUbB6AS0yOK/VaBo82BOyqjhTAm1v97SB+Eu6
mKpKsZWxX5WqSQq89aH+GGwetXHGAyIYsAgWbR0InDKE6ae5er3EEyXXVsgNC28GKlftl2Ja/fFT
PuoLCMc2QDFgaLOEtyj/Y7U100tnTuLGuGY7JWyw0EC4jhSoRC4ikTPwkZ+Lnq3/Fb/iDrPDYaPA
Susg1S0cVmzPAPc02ejcBcv1ccAYqOhIiwX+eke0HHW3fQqwj7tW54B94qtUOYU1lhDfqfdSGyJV
eJ3Hd/pvTW5XjtO7eLHohDWS/zdpKuyNkGrUvrnIWS6Lr7XQhkyk6VdLiY44aNWYerbMRvYqWkCd
7XFF4YnJ6Ej5PYS5AGfCOI9baGbTSJpxdJydM8YAbGDsE6IvPe4Tb98DkT8eG59PZb7672F7VDBp
HP6nXsMshxe1cmHdWl9je5xV1oHWX9eDqhsy+/aCcwdDnlyFomWuiJbbuK7BU1SbM8gRl18rzmmJ
6c06UC9uxafXD3gv08LeMLO4CJpgD9s0e/gkpHz5DS4GS6/QshxQE7GyXFepNGj+JD+XrWLW8uhv
1CHtdidzbdDTjEUkIHsiX/dieGbiJ/7ZOWZZgdOaswr+LMjj8Kw3gS0uTvRwUej7P2kmzLF3+195
TZo9ZhED0lfzXAlD0UqhAW2MOqzyP7XlRGye5AaxD7N6AaYZKqhVwky0ViMMMCN/FZ2yrHwMFGLJ
RSME9dCHYFp74D0nvRlzeMtVxy07IDUS5fKMmjK895UEPTV74HKVqQctxJBBeEpvvUkO4NmSL+Ok
sLhvcIQYso/Nx/8LSL9fThkZHfCSPTg7I0y2ECnlzI+J+olUDn2jLtPQ3j7B88+OAnku64rVFG44
EazTpzAxNVdgfb+g42gktfOKsXZ9yw8GP6UVdYct7xt01fNQc4HxBTVhP4HksAioQ+DJTi6ORDEV
AeaaCShgCe607mc30VfWWdkyzpJNiZkEbIsN43Lh/S+sCFPrVrMLpBM4BdpB5ca7mdJeEc/6+7kc
IVWs0fElM37MF4I8YrYWwVmVON2+aIXWPJOz/oDfTPHz5oYiTAnj8MsQzTq303IxAscAonskUR/i
r8VPq++wf7p2oqQKM3LTMpQYV2vGfjvt5E2qmqi2ApHgiZkK/7I8EBLyJQLi9fs+VEWHipxYNKf4
oCYiDrsRkDLP2/ZHBnTrHeX/0/VkNuhJGQ2w+7elBLMXzwr9nMrnvsSp/dkdtQJrTZzGKpZ96G3H
b7Us7BKsoYIsNhFiBufOdYxFIPbZzfGw/4zX2GhXtNb68baUdSVIkAP51a7EJ8XE9uCZccS9KQ6M
MU0L5Vdx+qQxtDBvxIJM8heGmTiCMaE+qc0ca0mO+ySrL+tFmQNJAm4YfU4hQJzJ9mqn6aKm0xRS
UTLXuBTHcrQufJnj/F9H3zPTjotX5JS6lyxrlzLZyF5uMr6aYIxi2XfRCxRffDL+homYdsbzEYMo
gIW2kCUtoKoAJviDCnTrd5NXoDcNRpkaZQL96eaWJNdG08EwZHQvZqGdqAMKXYgiXjk3j0JBGPdV
1I+FnPs2ydVbHFdrGxAT08PQEa1jknbiVX2jLQafYA/aVQXYhoaZxlgebZZMUu39wWmfqFy+jkvm
VRdJXJz5uXcOyJQbPkTpA2cddn/YxAtIE+zoMGEhsmq9co+3PsMQ+Qxn0+9FnDTcQG5jJ64IkteA
lCdU03SL8vnnIDLaiiX/fa4IoQBCK+HjZlGirOZh2aR6GfFKTwBE4TEULbCd7Cq+PM0M1ch+7aQc
wEycEgxgwJneG/1emNoH4xbSxXfWyUYYD5oVdl9VoZocPsoEvkKaTVCNIz0Iujb6ONkj/A6nknkF
yRIOHsU/xxRkJl+7lmMCHC/24ULxLOEwM5UDA7OGNxCF38bfOTFOPSVl9XpFuSnFgkVlxb6FS2Yk
AS7LsJs07/uAz7nDLbBtiT1086hbet+SiwQbwOkLSCcZebvF03jf2gALii+YUVJfIuSKW16zZ1D9
PvQMK1sH7iJORfq5qgJmuWvuQtBym2ZYmivuMzV8Yt5kpSoz/5AFr9tmZXJ6MxwR/dm54bnw2o54
LUeC2MFLMTBoF+xaHqyMqA6rkiej0q3OjzJDfZvhpoCpcsXBL7HnV3TLSu5DUMb4vlcJTbOJjLon
E1Bg1Z3mvt09kj2NErBIKb0sQ9jOtQ20aSYCHYOosrlDeFBaO2dbmYY5VONCWg1Ce46v42ZrrB6L
vn9/PP4gRmNLFUiL0KC37oHG2C3klQvlTSy0AoGFY7lL3tqyq/8ENFCUpqdg+vB4ZyRpC9tFrTQN
1jKYCgx6gkEVMMk0te2ZawbUc2O22MuZR4StWkjWJuiLsFhxroct9CIpTMvzJKY7YoffOOmwhHwl
xe1Zexg7UD9y9wR8+la/kgs3wsoXqZ6O/i91HchZ8Miw7b30EIWBrgvXbQKdd3NWRD3sU619pK+6
g9+6iwQKeve+Bz6BRqDwCeaIKQBfCmy0r0II6pNgvz+ev3Gb971PYqxIeUMuoV0hecdJ0q20pHaq
qTYT6uqJdYIwtRtV+6YwgZMdXemtYkp9Kz9DdLkTAfsu4NXjtEx4HmLRmkNLd81LcBr3bTodUoXO
F6f83bBKPDfbw4eOQyY+N3CcAU1Ka74qj5gepA2zVIUOOmXhv3bPhcnRPyY49xsnlVox3CTbmbvC
5FwUBBTUqUzSoiC/9cfcbtm7mMtXC/9Q2hfidpo/kTlm/Sc/GcWCJhxbVsaCz40RNTqfPEYvJ2Tz
9VCrLGndOxW+GJVv2UttQC2sDjbzPPOzVdcway2vJjOzg/9EhdMIiVoEbZQ5brlTEBcQo8T3kNdV
dr3mZHJa6OSd7deu+HE4KgESx4i/YpemhHWG/qvyYKO/oWw2w7q+GHKKPxJlHfxeUfvjDZgs1t4g
F+2ljWI1F8+nQXHYw7iHfx7pHyc5/Z8+6GeRWlXlSTDE26G4h0/gv2tjR1/pXf51COqXfN19nfVe
gM23YAP4H5s02iltlK1DjwvW0Cm1jP9IAgTFJiwlozd1Xz7SnG3ZcWP94TvDSk/++uK7lQSHG3r0
dLHkEizENBxadKLcXMQvjJ3YbKPRUIOSS6OpSLg+vnqGB8o2dHufZFD13PxKNukKz34gIRAEzhTa
v1Gyr5Y+cztTCL52+99Ecl4I6pp7i5o9D+7IMHEGKb/yx+GiyeTEM5GdGU62OdpVUyhjDChJwenA
/GO1A41biJe8JeA4iqgOpCtkCfFuK4Z3jQxInyZFqdwPW55xVJ5s8IDtTbk2RoICm/TLQ9k6Ncaq
c4DVydH0giguSZ75+X3zWzB01GspjslJK6YvrdJB9E+lBT3tIXEakM35U7G1mBC1ozzRo0n8JI5e
K4MP1zqVnL0JyO11IbpgQ8XGyLjbRU0Vd/7f3vVgcu6WiKiSOeci68QOHL3CfFwljWEP/BynccYt
s7mSs5SEG/5KcS26ilEL5JLzVzRDVoL4i0Uv/s41eP7Ucb+0VtB3pBu6A79L34G3Ln0eInoQgehY
7WeUUofG3qFLfZkqiEC32+YTym2cCaBTpr0xcyBQfqfGAOMzTYQdcqvab4syNHiRHcHS5gDRgCRf
FYjoXl3sSml+oRdpFwi6tQOKbebHFLF7OqfrVxtV4l/My1uG5VA/4Rhm5R0JdkKuIhsZ17LXqcjl
H/UbpQFh31tjfh4DmLc1iqWiKtArh7urAtp/kABZbUKpKjIYcavSA1ZthLmayBER0etoveuJwuhZ
FK1V8EiF8HB/oabMefv4gj+QFqf+yY85i9OpF8wy0C1HafRReU4+5c0O5ehNjB+YMuavklWXyRQs
gPpol66SIGJ/WTQwPSEBIV8NehA5k1AjLYr5ii5cuKFHC7unRZ8lvrps+Zmkkm69oL3Y7XDH5GQO
fssYclCz5nKnXdn057OHbD/4nfzbHAVCagi6tbFDcg1vullL7feaEjVC4RLxm19T57mASkGPYCny
KQ96tChsJxbHGzP2UgcwHTatA42qWXV5hStaOqi2/NQ+UVHiqvz/SVQG1TIVymSsqUA72WrOZQyJ
xV0hwYs7Sbis6U5pjSqhMukV3gvtyLQvXCvcjJkeXb8VbQo05ZKmKL92avm3WJw+PiEXeYH/i9Pz
pWhM8dy8QQrvuCm7fWFsOXHLXJjI6woZg7TovaABQuwTqmtDayfBs4b7j4icYL1E2KIsT9mlkXQP
6Q/5k51KV0rFUh4wXbesOdCPRuup2dr3LkuIm4ap5Yqs8cuTkzBXHfmUJShQSxMvf+UKujm87+Qt
yOxp0qhgTwGWOxeE+2bBtUXzC90Bw73+nN4Y7e6KXFAKueRInHw+MuDCqX6fHSjfWPoffcWHoGie
0w1GrCH2RnFsQnr629zHszWhA+Px871BRC3j6y67LVsbmiyo6AwJZcaLoaVlYVwC9zCJGkWJBGkn
xJ5tKNpmg3jQ53BW+Nbo9TIlUPz0pOLFO2fx2VZeWPODlk/ucXtm3YQIFhsg8fEnJ2ufTRR3Onc6
u8LrZicANh8OOxjCRVluCGuKIVl63LCE24eGxNNS1DHyLwaZ5FXPVZnaj0g/pV39kEdgmrARxgfa
qW11NpLda2wPOh8ONmUZio0nok5p1J+Ge8WfnJR1FYyy2qjS3K7mg+QnmqMHaj3gkX59wxA5oOnH
ewQVyoZFvjTLP5lUIxyeP/ZHxr2xno+8S8cLtKPQiMFA9TR8awqmVE9vIZ9TT1MZt5ksSMh+/aFf
rBmWLO5sBSU2tlUsviVhX5CkXPDjW026eaQLNggsjtSo7VaqlcPDTPy5NE1IuhbNAOx6ou5JutLp
WUcoMTux63x8zLZkQevLBVTcr69RSm7p4E+O9M0ajS2/PwSKwkB28pXNSL5tBpaae132jNJMIhWZ
ebFOenfhBYM7UknlMgPpEAFZNcfcJ0j2Sdr+kpyTc8WWtY6FoeQ9rop5vLffVJDqbc9n4s9J5Gpw
y9xeAr3BDnLLSGoHUm033zK6AXdvIY82imday3FJc9JWCLo9ZNOR9fb3u7DKcCtT3TSfwhIarg44
u5kZC16BsCFIl+xRryrRXXgnKHwsTzgy6EX/o3sZ/lqnoad2oW3GXOn5IeQCn3MGGHWvfUb011Rh
ZG91W22Mng/ADFuvLQoxTOfe8QHk1EKTEY4gYfD2KxnowKXHWdMRj2mP0HsJP9gE3nSArl9i0wdp
FYRXhJQQP7Svnk/MaqKnCK/tZcl3Yjwj9e1w2ngLEsf/4T77nivt+oqhWzLAD015PpAP1Ximytt1
AyJrs0IUdkwR9ExXOdZ5Kugr5zyitS+9XFd0zm/4rhFKfbh19sZJ7qfWZtEHY2Q4D660WyooZbSc
dmXP1yC8+dazi6T/qf49WTYRr8gxZTbgqVxzIG53B2wfizTwtgn6kxm8aorqUoyt/kSw8OHgNO4I
RGqj8wXBuIUuuQSUp64rVinMjz0jp8wQRbVWD71BqtpSrA2VpmG4SCuwi5Dbom6OziD8v4g8vjye
8PnAX2nGfN7spjsCl8t8UjuzPDnUg9C1GwUfbrraCdhie37JnarwCcBgDvnmhLe3iu5HDB8Tsbbh
l7TE8tqxre0ufKU0A7HI08dtfph9ec9/18qapRU7xPm7W36NeBHtKhQ0UDwTCxyaWrQmml6s522M
hsPi0cWlmqI6dyq7R5wLzT8dV+vdMTDbSNQd+w7evjquqK1IvWp1P82qpVsggYjh1garbUic5EeF
yJyZkcxblQevi3mCNjWVyHB8ds3MxTMc4nBsWvh6ns5RhQfHTREWJwKAbuo1GnTxOemU4CO3JFna
VeYd5+PlwA0KAMkrck7r5bwdM1oUIWlpx8c8ypqDVEr+tDXl1cBADfnIuWGXGKe0FeljjbKkInGA
9tAw24Mzjc7XfVHXNKKvwj/mdvzmd2ogx05ywmvmSsTskjRZPFiwORVCmlxmRH90lhUWveFdi9dB
EGduzxMupgacH22Z7y4UaAX+077lVmOLv9w4kvGHHPDAGa8YIjA3U+rVmEFhySZik3YpGbvg9QH9
v4Nhx4smUIVE0BGulzMlek3is601iMcfB59t4vDyZig+H613IC1Wr1PTBGCvpSBTkMSGU0dg8fD6
9N4rVqIuMtipW3eSCYdKu3FWi1EEQ1Mm8JGkttll7Wp1ISrXh6uNtn8SRmsqPE5ohsy/DO76VQXL
V1UldcLXKMd9iyocCyXLYf9S/joDLy7NPRyVX1Q9qH2Swivhrgb+sruGmH3Opt0F4O79skx0He4X
k7ne9gk7VEfkJP7bKO7STlE6aL8Jhx/kNLFjpYuOXWlGjY43cnid8Tdl37uxEN08uzdlKmU3qHSZ
s3FwhmuL2h5Mbp2ojbmno/SFhr3DVnFFnFfR6t6TeVqWO0td/WuCjHNsPHbQ7sawhU/5NCqGBG3+
pZN8uosdVFpIt47L577YdAzMGflI/pT9Ngm9BG/QomlRuqVhFdcA9+eRZ+ReQcjwseftiLzP3tYq
JFC87h94vLc+HLFBqlbbjgSwF6HmQ+Hk5F1TxO/M+F5sh+7mBbpCzZdVqcukV99ZG/G3wgV7uf0G
hWOZB9CLBVQdG/eLqEszht3+JdVEwZsFdJPTZS/RRluWpFEC8Xi3e3mux0dX7oCj7F33cqB4HuOG
JA+ftQ7jPLOCW4vTAZ0734PMNDxP/JntOonwv5hLOfCC1qaHu0CcvfAxxXDLHqvtHN4bNwDuEEeN
63suiYOqd68rKETvRLLc6Cc9N+TI1hrNpTmgBDNoSGUpRc0BY0BR6q6g+z8Y9hlHHFcLRG14d1K7
kJe95CQYD1war7D1L81CoKpoaxPa7TIipwsieJQx5/DPvcgJ5CY9piUiT3gaAB84sBB5xmQ4mMJb
Pvd8mdo6rx09xpcJeJS/BxUClCTuJ3BCEew4bJMADYtkcM1BTm+oD6oCmKsvKkaACS/tJg8JM4jO
iFlVCKaJyAiDyT8jbhXvE3X2I2CxT4b2fjT1acS7bi0UjRVYJrYnc5JWfrsbtqCC7+HzES8hc/dA
ZUGV9Pvh9J2ffzRbi3JPBUBLHAuvtVboBRIlq7phQsZNXcnzutX7XxtIc+tzdhsYwuviqkuZ3eoG
jEMF6H14N6WBWBeYUigza96gt3q/PlvqMdY1uH+6Il1Ckn7+T1aC7QolHrK2lohRY2AKDjU1JHFy
Anq2NwQi3CTxgaVk42DX8/8MCWsq0SRXbc9ILenyxAZ39/eP316B9i6Mp2wWx9YJ2e2z/ZnZp3Xw
2UhRss3cZvvIUaEdxmnhTtHsGQmJdHneDL1VJjCpDyRjQzora1aIILltxrG2sFt94nfCc6+8O+02
Dv14as/8ag8x8OowQ0Wi4G9LJkz7qkzNky1ZNTH2BvIfFoDce24yi9SFqOzPGi3B0rKoVn/PbkJQ
XUnjbpX08eC2vlsYhu5qaZAxH6nucqblDx8ni/mngqEG+vnwehRS2ztpoFJyoUC6j6uA5Lj64AO2
6WQCrgOL2E55bqTsx1wJF0+2Ft6If1rF8BRqkBdJEBqzNTQHMpilSMosKMAxL9ez1mr6rTgvOIye
4h1kVMQlGiPo7HV+J7G3Nz0QOUp4zADQMM3IZCIOkbm3HIah5WbcVVcixADBMv+crTnU9uGgtEKp
iXVLsg72yPmqIUNXLH686DXrJXSV+BwWiurVVjemBg7n1Z3RoQImHrqGy+o8heXMnEDTPrACCXWm
LZc8Ui0dQMaAMYXG2xtMHfDsBTQRQSihJtE2xaTVPbToJETs/Pgn9lfWkvuVb7opU4lo4LO8VPJD
kgjB1ohOBqRXZ+O+GaBNB1Jm0YXr2xm261W+ezJwSo+l1CvBAnC0U3K99rznVpKLSHOsw0ZlYPlt
2/FIqfVY09afft32nEDeDT4s1VerNovdZ6T5Q9D03xq95qBdcUeYSSToAtAREBnUMIV3q6HN0jTX
m0o7DOTdzmhGAdA4Rt07GsXRCPviL8OJaINHtVmuuO9M2QuYu1a48BgHBB0fYaj3PUdaduAxVEd2
/YqV3QIqKVQVbuEJKysV+aO38l+vSMo3QXV/ItnzuMu66Dd2Rpv4w7oBYRpM85mB3WcTRgNqD6+K
QMemv26yJ+h9fSD5Ie+JqDaWlDxupbk+KnKrRl+y9nvQUYQXD6ORqv4NVp7JS16CxC7MG3VAl9wc
p8qo2DvhXxZ03/ahaugmxeIprdoIG1bh9xsncgIxXMoJP90ic0d+0+DHLysvj9BHIkGnAGPx7CgS
dDED+e5al1tqMbqmtDxCapnp+oO3FLIIbKdXxtcGhnjWp9BOB46sRrJXad4etQ4ctxEFye06xiWW
jAhQuOpe1S9yEBaMn6tDxLTrScYil8QYzdP7exnm/RNoN5/VXwt34tkf5D7yOz3hmlfu7AnNE75y
5idqAo0o90Af0ahMfHQ10uBgZTLlB0Xo8i4aB9d3u95ppcNoCw0kJdk/9SvS4OKR9R5wVJuTGk/J
xz5Y1Hy00Pcu+VRlj0QLqRHmsNhqqO1S7RTYqXThXABvfki6rkNYC/hpqqq0JVLGVJLOBmNkfWxF
5puePtu6ey6KD9Y10U26kadGFPA9fPFc2h2ElkArJCI74wkfRTI1L4NooL13bOKPdqM6l0XjQFQk
/lxLfjMCmZqSBkH2mgChSSZ3fToKrobTj/KkpkUA8VPfGi/AyltglxHE7IxnM4rHVbVgRGuxAWJ0
xQRT6BMZGrIzt/d15yuDiYBbpmiBLzKUBJj2hDLVZgR2iHzMeBBGl+tqiwrGIjUge+ded/F187eB
3gvR6Tka305CUGAq4rpJWahqDHEGBCPsjhoIOz3SMJuxYTh5J7WILfHya2WVGvehLVlM6joYqmn6
guqeGkEsEntndd0rUjS8wF2QrzKMBrdSbv57B5hgnyw2gk/amorjSbkhw6WXFMVxCRlDK08Wluso
K/B+l51dUXrXMqauaPGY3IucpRCAk3VH9qxGBF6qV+7HlsVCZMFLfo+uQlbaOxxGcYjs2YxseMYU
8heV2P+132w5w7tyvy38cYgLOEb0jqy59ViIOZyYSlMCAj8GByWi8FktbQVCv2Yycwey0UoYDJ5f
o27Y4XwflDx+TtWXXZHXqJJ9AYR++N8uBA/9T0u3n0yHpV53GKSo77bOhud99KhsJBpxyVFhLrEU
cOFYNLMEaUOAaaHdX50vlUWz7wwp4IDnp/BNGx72f2ESzTGwEnkEQ7e2KkYiTzHqdONK3ISZ48LJ
K1OUs1cZZO03ten7IJrx8aSvv/mjj7hHDr3p3Wn/xVW8jyN+ggKfvjH8EZyhhtgMmywNsD5K+eg7
HRkZK/J/mKaQ9MC9vyV2kJMmVwHTwjtog40dCgo+mMgXR/KueL+4sDuHJRWd2exskTnjf/URfMsy
vIL9Ptl6MbpD7JmCO2E6/6LqZuMf9iP3EpQDZ0J7/CNGkausI7g35eDwNXno8OmlCEQxVv5xqL3k
50dB4koeHBv6XhMdiECc0MgoFwDwgY7ZfIA1KyV6hwYNz/jKSqFKZb3B+ebPwhTb2KVhjLzlZC0C
ibqAzzi9arFmz+9omyoQAiyHNvqqhJv+iMpbCZzGZHI4peAoyUBCruwthjzt8M9nTOWXmbgsBMae
0JNnIlS7utzoIeC35bN6RrRKH09wcK/ceR/8AHWzcxYJ5Ho80Q5442izkFJFjnut32wubaTA7hp+
LLPBW0Azq/v06iZBhHuevMQbpR/9IZolE0YMeUr1z8snnu083Ggkkf9fakg0jOktOmZ3x2ytKzjw
m12wsYx9okD8I+Jh6J0tjKEIZ4gV5M4AR4csqG1tuTaxyClgvqfZ6MBODEjG0600mrTMTzwYZPuj
8bFO+QLQMeX9ZrARZLPG79xIGhu5zOPji58mblUu8jYwQ8mcdFRwrhvfwx2yDMgAQGGAUfT7YU4K
LhtcX8AsZQ37VIL5PN5ntpWrL7TRihah6Dx1lG8nxMWgASzPfWRr5w8OTBVPst3I378POVFPBPjr
K7tkj9hwMUxmi8RXfnPewptUFZMPeJV/QO8LEbRfy4hpaDXi6Wncy2mNv65pC0PrOCtR4o/tycQo
IDijNKx7czHJ4qBMbWvtEWH4xD6fCF6prrnB53e1uM7+7RkFsFl+Vd5izApX2EJ5ZbGOLr//W7Xr
I5zlg6YLuD8Z+Tt42DAiEc5apJwP8c1JVsIBLy+oOFy94/jj6QK+DOvz+kdX2Ihj4pkOA0zFDSrS
U6C1zCul76kqcwEhngUu2sujy9o7yGhVyaEa5q2KsQdcKf5mkSDM1Lnt9FMPuPy7/H1mqn3tQhKi
G7GzAlbg0g+i4yQylXH2jobs61ygg7L1C20oJtCJ7rijQqVLrjqAEeXFlEuQI9ZSn6+FUGD6L388
d0QK3+lneN0OCTjeDjMiOCKsbBTNOBDqiDIc9gDUxwwhPMYOrWVEdMgPyrWzIqGI5tVPGSrBpWV9
zU/NEUWaq9fKWagd+p3bBj384jMlV30wYMCf5Lv9tJy+mZpR4oqjrztWjVrI/vX14J7DuXOofdG3
4Gv7pDgs04goqZauprEMIvqgWil+diVFFbhgUy3M9662yWz6P1BLds7ld5EQYXDmAhzvrx82DV+3
LqPlmG77+zNelMrZ5xMhWgsiRmXGL5V/BBrmfdAnVxU6OZUg5kVCQs6IhhdbLUWCEgr9TqexcLRw
/BMlKZBsyIOVVbTIDsotyVUeeBUwWh/wOe6euUnpM7w/UG5E/5V2h9NckEv5TVxIie97/i8ds1oq
M6WdwsadAjm8ltbPwSkdKOAJDGl8U7DGGbRRQ/ASRYieC+fGoIk7riVYQ0HV8PCX/fEfHp+ObLD5
p8+E1MugJhoS8eRa4MmTQ4BnEH9GBVzAtqAbtpUrp6TM6K73dqYEuCo50JjESLfPbaN461AlvYfF
LYwQRHedk8q42dK67ZlVBQdfL7zE9f+lbzvU0xx6AbdW5/AgQf+SQHAZNfSUmfRKduPCv1VmXpND
94fSuyTJm9QLrY3Z2Q9Gu9H0sTLXDVo1ypHjlh/Ba7pMDN8gx/YPid9oOtR/SiKF/lt3ghdT/pCt
/D3nbPzoztRCbClIIN0nNmNBp/jTmvd69s0IwkNVHzsFaI2RRO+VWi1Jt9u4fKSHu3qaXpFZIgvj
RLh4xwwNoLbCk8XsS4EVPAkz35ZfpMCP+E+lA4iaVN35UdLb4IsQu/3EGw9VwDpHHsBn1k48RLlO
505bNRDPrsznRSsbVZ9c5MrYUR6i91cYMk9D6C81oVvrRYSD105M+1yKbwnn4NBpCKPiwUi1ztnE
3cjzqftBp+G2/sBhPEtUm6EsMOtUe32TdRLL2E7SXmpeyd1VzWXetkZRQ0q8XXIRS/EgSx0xKwHo
IG9khi0khI0lnIXUO74FZkj6nKVZBuqu9knb7RDGPmeberm3AbqnbyTqD4ETSADbYmDhoA3ilnWM
c5RUtnsf1SVMQR2RBiuLHQ66UeZjp/gHcTTdlHiMnFdIlPGHsv1A0QPEqYlFVpcNaDzxoqir+WR4
DSbCdwoMGNYE9mOCkGTFWDTr2FTPhvfM3NtbKCcpFn9vUuZ1pA9Lcr94GuSlTrGKUXI3lyyoC3bW
oHbS8KvN3NsIDD/Rm5jZVAqi1yQff6bGhRBMKywaraVLIhaMgGQFMxZtqW1x49J+APIUZWGnM8yi
WHbo59VnHAk0jCiY4AAGbUl44anVqXj+lGC9SB5ze2qB84aFdBYkiBId2qk9YIgPK88j3QPlqL6l
ugt6xo69riNkhYXO/Y6mCkH5Dwf3An28Oe4mgqGGxLF5bEKRGYhFDUx8Dt7DsRWiroyXlqMj8tAc
7SmonDuOuLSYd26+A9Me9l8WFLacknRrzoyAC6a1ShxhvSw/RsCqIWh2FAwS7IG77W0sdl2nbMd2
XuL/bTY3EMcwaAJGQRJ9i7TegBpwoI09lhqZba5FA3IzDkWZL5exw9bg4bYitOq8w7H2r0jPhtdJ
9RQzqLIhvU4+sdozGtkctxRtLZ6nna3/dl8TTLfRmKuoByMbNw7hcdzjGW3rHEBA8lSlzOUfTcTj
EBaStJWpWAYdFGNHUqly3ZiBZhjOs6T8bRlKnbhU9wm/uVuxbDkq1BUlctnCXFQUu1mc/crTo6wS
yNPVy8ask4VErGQ3xu9rumwZspRwhtARvtTTPJb/o3GCdcfv2xw8cMeW/E9zOwz3gNJo31nYnpkD
ko83YNiFwZny2tJWuBENgK/j5X5t51tHmj1LLyAuBTi4rLm8FpLFz7hM5P6se0wpJkmBgzcAmcCF
PuQqzui15RXFCkiyVKlmLx0jMlR7AUhwN9XSAYqXKDmWlFmOpnyaSBzqZyKgPLkpdsCVUrqpdLXe
JH3kaQRuKFi8A45BrcytL4LGUxJPYMXlzUX7Wcop/eZ9byXhGM/fvlLimBWn4SapVAIo9luKP0BP
iLCPsGPIVXxX0mmK2jvRNqLQIiB+S46WE83b3tD5WKJtdQBzvH16/13+A7PitQHIGxcyw90Oo32i
Mqrg/F2/xocFLmOyRiWJEXBXCZ+0DFVqg3Z51/DXm40911LIySNvIevgw5DV7qFsCFGA+sLkfc5S
AH/R41dYolrwZ6nZMhWH6dtx3CI5n9KoRI2lFVXsnuAb/8uPGqPqmq8EVKusz/19ZG6EnQiimBo9
Hd+lq+qDS0etOAGFuuuuta0dAZt+y6BAoeliBaFHTgNhiJKdDeiVp66527X1R4IvN825gFGd2Stb
5bbMbglKLFmDY4yrncFtvDaQLV/bjjunCbfVYI+IcrlXlTV9IQBmHwPstzYFKDpqzEWwwrblPnGw
1Wuy4S7s/0wz0bmPXrZyRNgZCKlqpGJIGZTk5cELnebTAI/oCMwfXM8AFzTxSgpx+Zw61zVu3PHo
VUcLaXgA+VyVQfRqp2t813QpThVOi93m1LOCe03D+Txdqqdbvpss9gKAr2Es72QAud/UUxnxutXv
nzezTSasyPmMMaUYkvZ4P1Afe6JRAFlkDyJnTR9ghJBwVXOsxIxTxk8Wzd+U+3s/ou84XTy7UMEK
ysD/JLEmFp3vGvxBsKWe3zPkWLjZnhzw5mxAf3U92mBIw6EP8EKJjjn5DHtuM+pf1NWiGksQ7DGf
9jQlPgWbCY8Z+n7jYMnSsNqbeteAhi9NhHSdlvZPVHFr37JNvuU/vQSJTLG3pzLBfRVi0vM4RYRJ
Zi/kFL3U2MNglQeC21HjaxvryGrJ7fML8eSvWA8VBv2qeJzUUQgyEzbvnOSr/pGqrJOiMTCL6wkd
cf1Yqvyp2pIbhDoB0vQTWkRA4ZJuwNWXLJnFi6GMeyKmkuVfITE82nkPujWD9Z4nV5cEHuwjCOcx
f7BTwWwW/5UmgcxgUt+YRv8XT0jounQlo3faM/jskQmFvQaWSYY2rofrHz5jtqKPQH/RrXqwFy6Q
484xHnnP27BrrmH6Jp2bITemVKVXucrbZ+ibea69hAp+jok/nlGM3UoXj4L7vXJxHXRs5hlCNiLa
gcFnsV7GSI8FwyUIyLmXS/pKSjTMPPgOTWYcV1CpojR3POaufn/EZYvO5BRTEt7Ds9HQikj/BVcY
DE2EHgQXnXOVHhLtKiOq6h57y6C8lNXY0FmF9dMFU9LMw87v+Bgf3mGhmHTphGMaIlZlUzQNhHAS
h6wjXjdvQnzo7g6zkvfWyR6W0/8hHwIk9wOn2nv36D02QIA+ZuMzfbJv6mZN93lHXb85eX8MBx1p
wBILgFQv9wGupAb99vqdePrpO75xWcNp0WZLbk85QapFoC3S2m1UYEcWyMpXTrElL/ZZkwIIh8gy
jDYcujrIRqgTSANCU0xNmHAi7NE3d6t48cB/cSm/gCPcaZViO9r2tCgtPpdA+FN6BWeXbNBOs2g2
15vYKMa8PHYeD7EIE/65MjHyI/yznhylMZRHZvZQl6HTp2ZoKtsbd5dMOvVZHOk8k6Ygii825w1z
JXyaJlF/2CU5/d6ADxbR2BwrFcdXX7AZGQU3AES6flZdHpcD0gr0lnKRrI2bYik/uedN5HtnR43v
U044dJIpCVn9w9Z4aMJM/doxvIMwXYgAxKGe/XBik+3WJhgEu4CVCjeKo8KMghvt3X/enknqEN/M
w8gYC6fyOcnWCrTv4yLf+Hxc6S7yDzFYWDcxffV3dyOKRQabgSxpoLmz4gzsbfioRrewBkp+y6h9
rIYFOfngzlNO6dvH6ZwjiGbuZapv9+TgAzqEpT0prYkAMiLc9iDjl5mb1gZ5GLt/af/3T1O5YIc6
6T/+pkcd5hnTAJv+l9gp+iWfdprRD2mAiT3JUysh4QF0c1yIHRQ5ZDTPE5+4wknn/GErAKL74kYt
bOxMZIT/qGxlSc0i1R7cJ3PxGycJO4lGxC2oJeGRBAEIVELNjc/0sUDqMsMhxrbMQ8kwjIcJwVc8
PhcBrNTFV9dUX30zaITr947JGy0GioJb8mKcYvARcNc01dQCRe2QlWuPMj9fuBCzUYwSsg7j0daH
Xc2MYw86Of4F9O7Ab3MQaldYXJyIiJ+LZ+rjN5WbDXvbvlEwSAKLPINOrVH3SsPIy3YMkxX7X728
8RXY8yrxXvauGAVKhmTZH9gYe7x5PSAOZ1Wg7GTJ5prW5mYfA56DXplccyLMORxaCHAoN+igmQIT
qtl2x6dQkPlALCVGxi3bcdYa4fuKp4/tNed5uW4lZzOzfuQb4AZJgrVt6SpTYsHKju6UteXB2enW
OG57nCwWmXa2uXdf1sHc7ZwPvxxXuE8f7cP5IPwFSMBFLDRvuYzi8DCfn4MvQEu0SyRJK4/U/Ljw
M9ehbG0jLsbo6cUGXu7DKQ9n1PzW/CXnI68wHwmSGxQb/DI2AMnfaKCjdQKKGFyIKcdlXfPwDckx
DfxlE2/z4mjJwvQDUwHhbWIeCyR1xDiKKduFLZCxoQ==
`protect end_protected
