`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
qqCrkr1tFvJyLhqq/RMWaxVbPUY9huaUkHXQJUcqf+Sg2PTWjMFpJJCyLQ3N52wocu85IItMaA18
MhiDs8+sWg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
QFZSghpnHMJqyCF3QvPSr7uGnGjg0heEkHAQv7qOQ43Af102z7EuhBRNr64oIxLGqyaGKli0g3BJ
QkHnKyzQHLfmgiYU3rxH4QdDOXW9R4bzWQPVQQyyW+DRDou8+17XFqq/KJ0LO7qFH/sm+AMf0rFQ
//4AvNVUXwz1lNoFs4Q=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
wZzwMHG7xDj3H8aKkUNc/WKlqvMmIxHg8sQanfq7D9gJkSONXMBIO6pPO87AIGYzLvAYZKajqCLH
GPHCOMvf6N8/YjZhUrnxHhRD7jRRQWUeGSD/FAy3wAlzD5SQYw5BN/UbdSYmRVoeWrUbjDBP4cyK
jvwxg1Q8zr0uFbdyQTg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Yc2lnyrj1dy1fM0GniWiVc1ocHufSlcpbPf1ZUuNv8SNOOoqjVzGzZ1oD+Hu5ZaCsypQAx3o/6MQ
C2FCJNZOTzj1fwgp2Z39ST7SeKnvROX53Gy1Lceo+gGr6z47UrM2LNvmU6+UgS4XKZNhX2q3W2vg
2dWJpZ4myQEsmZMvdbx0UeSJPYl+KCLBbrpekvhzv1Ag1SePGSRA/tV6s7TMNNxM7LFykZNO/saD
2jL9MgQ7Qgps8glbAr/C5d6LYpiQMhY/FoxCecc7GDwYUdht5uqPQkppiIZ0cILF4zHW2KvN4tqc
4rFUMr12WjQ4lxKt9ud6jEgtZNq7i/KPuY6c/g==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
hSTuz6zbMVD3JOZezaRgjNt1UWhYCvvIDpEqYzxjcZ3bTIOlGSKpfCDYXVbNvqgxVC/4Du51J1IO
M1gPI3tYurwGpYFUlUU/52zGRc1VSOVhoX/Wtr0jpCZR2EmE1M40FNknf/1ayKkNCSOMcx8O5zb1
lYcK5Af43lFrBBiDiWH3x0EbchTAqD29KJfcIP75glGKJYggSj2V1q39K9Pfs7ELG+LSaSOiAr1W
k5Y+ZGnvmzKJrt5vyQ7LSG+7keICQHvvh6UUiNTEEmD7Fmj/HQPLU9P9gOgdYP5XI8wV51PA3w1Y
bIZpMPywZuLeJ/7MTuwdiQgwUs4Lw5jhh3a7xQ==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
O79UmbhWfeqh2iRYouu3ubiaRla891IBPc7gVoNREY7Xr1FjvTzkj5QPnLZN1D7y2ikzBWs5Qif2
HlYqjWGtXnwAHYXz+SwqDtPm5YwkX5VotPEm+AoM4AbHONhdQ2SjSOWX/lX9FHT53wrozdiDEZmd
rffUgen1drM+ZdmE76HH2jEC55ZUxOcWlMtrwFSGQck2RnJJXHiodhzt3gf+FbkynqONbayEJq+e
z+MNSep7vinDgErkRnhVuB72N88LJr2c6endKeKZN7lEhFsGfFZZ6DgZXMAoX6L2hMDN9+vSmPfp
2M3HLgtNpEA+J4j5nVNEIx8P1VPr9FTafi+E3Q==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 22944)
`protect data_block
FUUfLSVKK2+6gSTso0V5c5FS8gBFyGGkRIJuM6Au97yiPOlBjqf+M8LYZHZG4I0QkIWt1mvjzAoM
tm9TsqfwrVXbBPjOegQ8yGGZLybSEroXAlTtwRn4FSQSwMrNMsCLGaJkdAiCM2eN2fB9GXmNWg6I
myr72+HaVc6xzXV1VZPDn+Z3KRX/7TnfWIyjfbvhZkr1nsdN4tP2BTXbbq+Qt0zTAlN02nPQZ5EJ
TMXiItLq+UX+cZNWBmsTmZaZagl53a+B/EMhwnIymnKKWEFWOhgnIAOn/w27RH+zFRHdYHHaZj0K
0v/zSYvGG90JD0EcQ9DH0COtWtjiqr3rgGFIWxZWls7Fa0Qn9U6cSmH1A5nmj2dp6Q/9e28y4ujh
8l/hfGA86xnodXOrsMf0jFkztASArvSwmE8/e+YNWYC2J7kfokduDZOSdW5M6vkWTaJ47pSocKJy
Y9gAsrWe/73a6YUEePtBYX6AY0+wDMM9Hgg5JHME2Jwf5lDhSOA97dmm8KIC6JSv3lBlUULhh2et
gzv8SZSjRT1QkBi8qRGc6qTUj7MuJgD1R8szyLfIp8VnoA53DFO9SctV7LUDRaTsfvnDALEmszCa
O0uiGUfulBb+9jgx/XDbrIqAs26EUZtoXw0EX0LeuYVMVEOigWHLgDrfFbRMOxakKkw7Sui7ijYH
3O58/cdsiElKUIpxDVOu4vTT7Iv5ehGUDqQYzFcRG89sPJeRreHII8NHvHHVafTFanq2g6W/WeGh
Zan6tqH4GtYJdzHeZTnp3c3YNd0jgJtVpNnrt9Bf6WoZOvDiMj/5vy2n++p4CwqP7/Ur2V75GW6u
O7K2Yy1mPtL4XAbdbBXbODPUyXJZitJT+zDP8UlWOsiW3o/Y1WjQ3M/yJ1XWUCJByIQEd5AuOwfi
/JCwxyHwQN3aGNh+/y07DI3pubjxJMRIDn8jPe1MgBBN/iwe0wwD0lbcT9IJ/YDTLhRiIvaOWi47
dCNCbSll5KkGTCUhA90Yq2YuTXk+1lnGVLf4EJU+8CC3wnNRmQjX7x+iMaG3ykZ8Xe0f8yxiiYqi
henCTECdlpb/u4VMMd6mTu2D94lW4tqwrFKb+RuIpxSC9kIqDyEKzxiCiesJoDm03/llktdU0tJG
wrE96GCIQg/wghR/N/6W5r6UxMlHwOspKWbmMQO1qK5uH+or56f0NVS6E9zPrvIxVuD8shpOoi/Z
kM88H8sCcARx/8kSNRQZwMr9EDDaqssm585VT/slHmLaQm52cxqtys06fLhOxCdPWUgekE28PYgl
3uSVwete+Ek61FnXU0T1wcCYZ0G0SHa2BQeiE4u+ODwVQtC7EdQ3pr/nu/ha2qyNASTQoeewyWtA
nN/ETG3nrwEw6dn+QQI8GcDznILAAxNxKyz4CmwEzAfVYQQI8DQ/9Ej2auqJB7eWT2Xq0vyK5hlJ
ag+mQYrl9TRTcvEvS6jkkuiNAaZKxP2QHL1bhk2wmJydK30LKFVYPo+0FFjCjneKzYMgWGM8yLMX
n/C0ZlmF3xHwG4zboGtLdR9sMp3uz0w6+HhT0UWIWxlvst7v6lkgaN9k+kwJss4rLu4eagvAdv2g
Kc3QCaxM5Ne3RAMIGyHgy9wJd2ZHobTmtuMJt8KAy/yToJOxHEr5c0aWQu1kWDn88cM24/Ixw/qG
jAytoATnPj/E4zTnzDmE8IxHpk/F5o8KdNfoIJ7O58xOJEOS/09C/Sipk5mnXM7O+yhypEq1JCzM
RZJ8Vl4Uwu2uifqtRov5toVWfpHNol3v9xI77/hpUR5dDxIQNKsFchVfk7ntIo5CZTsYlH34ZK1p
2q58ct2GC2vWzjY8u+j8rVMl0oY1UUH7JtWaiKuppAdGag59K/pB1sQVSXoBQEoT7uEG/ooeJJ3n
WZ+YEMH2WfT8bOeKIZsUlVFIdJ5D5Ct2y1lkg1FbHf+ADKBdiD3TH515Xvg3DaJtNRMlREc1KGf9
i0KKtKIi4QEhf+0tC0rIXNsqwwIuxeIfyZgSUL/0G3k/QsqhbfVZOHncNc1Zgvi3VEbEvQdcjMEq
MlBUImdpN850F86vXrlzSXpzSWn5WNR1N9Azhuc8r4+T9/GoNt+8BgSATOffsLHBYnBeUMUkBP2B
utO3ng/ZJcFzo9VDNRq8hwURlChAPnw2+CUFjKrwMxKQet564gB34lG0gmoRTTzNXzeIwWmhy6BZ
l+ROYkXF5TUR1E/5qOGeyMt6+KkVGdEoAd7o+e/HGRtDVSAjd1KfIuPg4KyFwS1BWgqNpNGSAgEP
cg03k3CO4FM9Yz4704Vwgx5Cx4ATIpOVbbtyzSrD1LgS5w/21Lgge4e5QANvXh+myP8c3+2sb9gL
43tgZHnu5ybC/Zudwt9GP7JScWB1lvrjO31iEg7eEXU3x33Wkt/EwqItUxpVlSFTo6/35kByq/I8
dNbs0Fo59Zyto80fD85/Fc5DwfT/EiNcRaiVWuk4hViCd1G4DBsRgs1W8VytvAi8Z/bnMvbJjSuN
qwqfSJTUIrHllAAhjgcJnVmqLxYl2dOgJLtPSmblotH5uSHUACF7UR1xLcXBm0sFs4t7outg/KFX
X+E0stQkjk0f0gCOR1j/fdmF3plx1ENJQOcgJRE4ZiAIHS2mG+fW2fic0mjkxwwOO9wEinSLX71p
4tqNmj6xxnKYVuer7dkhgTOrKyxfXpSxFy4zhrCEsGASbJsdCe2eK6VKj6cukSFkqjApW/QHBubf
rRDdoTD4ffMiQu7Olj7lZUYgFuAyjHyNQVOjwpAjx2+ATPcPHO8fdxzv/RgTN3xPYMoINvcrXcIN
Llyk9OK1LcF2AImfeVxBg4ueap5XerWb6xlzH/JErXfBI1JW8wIF6eGZqLl9tF5rJIBfn9RPVWmK
0cl2LE2Nm3eIwfc1RuOGJhYUUsfIYhsXgFtZLSlTEWpe3nW7ABPuzrVEoXrIh+YmEToEKpf5yeZf
hu374l7px2znIMd0gHczqIWveaDiFLiJJV9jHvf8q8VnZUS5NODmhFj4vSfRZzbGKiKbvXlUHnO9
DtZcC+qpnY0/c8EASY2gLhd8/RjPOVHVdX6HpUdpe6xi0P2Z71abOuYWlxHYwqDGchRzA4i995/Q
RLWZQ2vL5YYn3fzL73LtDN0hICz+IPLs9tvNt2153CMGDBiGdVYzYgRrZhWHjfkaMX+u8qF15WgV
crgsqW1CRiNG1XjHsWReak4Xmi9+DcI2tuK8y1WXW0Dy/HXj47SF3B2b75ZzVHuU8SmFY0uW5RMz
qS+/bYdMiJP5nS4lyaCR0DaTlZDwjzuNLq7VyVkQIdZth357ehUq2eyLepR6jDEMhO36DqVEQdsT
TiQUAh9z/nulZRVhhSjbxaeSr9ATBK46BUNRJe6YQO2qHqr6mpgpcmFUgKV2rKn02Q3s4UkXigMG
IEsisFrLoJzsyIH5rSDajS3tUEz1kOD6HA4lS0aNB2v4kI2hsRbvlfqqgVwvbLapp9KgMsE4PXE/
2SMWEnSmY/donbYdvk8U8dibUkau7Sy/a5QzLBlMRdqWG3Iqvk0rJgzKyUDUXVisgeCojHprJbm4
W8T40jvm9aUru0SN7yWTlIkRFCnrvnSjuOJpZKtMXjsKAKvnjkSeRgHQQcjBZ6kNDXSVQ7/C8mYQ
WIi98NUSXP9X3ZBEjg7qZNq9mnn5Vviai+Ulp5hQYtAoUtr7Bic2OSMWa6Syh/w0CGcZ812Jdj6H
PLxR8z4RfKk4VI4kYYcNPUowW/fTr63n2x4oPha3UtjZdGZJol43MHWmckPDQp/PjgvM706uwKF0
k6Ad784ANcDP7diTkcbLXoq/0qv+yXfKL7QaTpMZxrCb9Mg9OwHbQWGJRgNi/QbMRad+XGTelyys
UBL+K61A2sW0nWC8YSMaul7tKvey8sM6tOvV9efMO+FtAPbnAwEYQJ8ClPSaVzqKCLgGgv1G/s4t
bz/8MtAVufSzmNTKwsqTg5ah+Oxj+ePzcwYetiM0d4OesRYu7Z15QUCFkl8FMnjAmoMtjiyBWHPj
i2SFOrghopTIG/IOgETcRe/Pajgqhbs/SCEUtf3VhwBAlaZonL+7ZeRSDc5sd1/J5OZe3S1FAAru
WXfhaKy4NAnFXjv5ZXBNmOZvXluU4vm8uXbZteHLtll4Xcw4NbfIQAO8b/0vz4/N9929XIoTQA28
s6O+UL8EACk/QQOsUfh7Eet+v42f58k+//9ejJjH/mbaWiVYXPylaqkNMXG5W5HYdw+a+Rw+m9UU
hjK8gL7glt4jkXmFifpSHzla962TEQ+lcuEeE+njcX7FFctzJWX/ctayfkRkvayzi/y+bppPbe0s
xkTx8uyuIG0fCSzGiq0ha8RJk77BD2on4rwUGjO87WLOGlWBJ+vdVgar6zugXqfIr8mDI+CnXOWW
1LeBzhZtU8ALK4ToPLIGwmjr45lE+S4dYfq2L99z4x2wtGXOnCGfoXneQ5mgGWS6AGIy8j2eneB/
teVKomFeFd+sOmnHRX1fRGGPdhyp3I9xRzCzCHVSNG4+ts3xClegEO7rkUoKK9G1n23giNesbEt3
FcMldGq683UizVV2R3aTF50aK6fFgiA5Erglb8vkzkylAvV+Q12uDV0TGgk5UvlCdh70G284X5q1
vVRKfLF35iWnEiN/7yB+H7M5JJdKARTdwG/KZy+nvovIgJQ6hlXyMn5rv/3JJ8UgpN9Nd6qtpjPr
sHBBcnqyfwQvotEpgrk3Rs2pbSXe+PrPPd23ZYtBO/AziWfo1Cb9FXsk/vByHBV87Fi9X8AjLjwE
TelfA41PjGiyLx2ZQQ4igAB3FsWE3FEimrbHic8X1pY0IhcJp+RzVJz4I3iNmuw24oFBRw/5dLrQ
4mkVB+B9GUv6sH8bYT00+1NDK14el9OwkWWmdBMVIgel1PpGhm1snYD1llw2OkM90vsRc9Sx4bv/
emTiFEibSg1JgUQVHp1BknU1VqhuDEl+hw8Rcw6bD8nqZms+UZct9QjvWCzQTIpabehPlLogqTXT
nNEYWP480Kj2RFKDLEjClD/RLrPHcCBw6RjMtrMODN+6EChrXx/nfsqWkgn7Y1FhFdFdIXiTYHnU
VeaFkyGqAVX1e9Pds/cnLb5H9RPZWza1y1GRuvQcPUb0EpRbgBakCU8kVoL0ZwcdVIeH+fCU4uzK
qc91jmOfViqydrC5uBe4B29fuiNOoildLW5GuobmmfxEIwiYA7lzd1km/M4Wx70TRrQW4ktS3xV5
RPWqbU5chLo/zcnUXQzjIJ4vt7t80rh6d8/LkI5v7XsmTJNVEmv6esO/m0jMiLsb5o+YNR5GnJTw
imvN2AjURCOW2nJYr2JyVjJLRstyOTire0bJVR3Y2tsUnziDDwEGGb7P4kmDdYOFVMwyb5jcEuzn
6kUvDcn3TQFoH3ZPoT5RlfXyyE/azsKPvwwdDJaFzkwg42bDukqp5vmYC+EnioazOhbPNc/VYj0b
2bV/1IKZV9o2Gq8rF3y605RIjCyHS5z/yVpbn3MROMywUMSXFSZsl4E8YZfnUKv59It0jVl+XJBG
rUG8cKEEzTb8xGFBQq1WtKYi+eEk2rOW8+8+UNAlWiq+25x9inuaRFAJpN07D9iknD5STwZajA6+
WlGQ5oCjwS37GWLFcsZzY1s/JkRObXd2yx0Tf7oeCynSAg2vbZadNZEd8Kw+G6BMZJzfgranhp6z
cE6Sv+3uzvYzYrjk4dljxpvcAa+2oty8UcFLbpjdTmJLqJxV4fYVhDWdqn9f6wpkhZVIZh26dzZ2
gWc6dsMV0zAZTyaIBDvA1IXx2gsFeDMFOC/5E/OAD6WviFE0Sk37cxi496thVKtxC5hZQuPkXmoE
UXvRN3N9+KnQpc5ZyXiFYsJGtuA6TLXQjbI2sI0qGPzKvxfSWcUW4SJDTjHgrz1HTIPHJFdifDig
0cGpZnfNL9b2L/lbk5BBMgSR4P9fB9jh+vsTWfA8a5lumJBHBAN+wwzaGYrj56rMQNuICIlVpwhb
y4ftJm1+ruJMXtVJMuwhF5qLL8qa9YDxLPgf0fLrVTwHhW47UTl7zBL2C3zqgMoDxbUu6lZVbNOT
t6J0D5w+GXqfRrfVS8mQ3owwyd3GPvx7YfJBpwe3lVM8kkgZmlLTzUq4eeCvhRhuul5DO20XK8ZT
3F8UWo8AOFTElESSJmN/2UdtmsvMVGTUTtbvo9e6HmcAex8yvK/KOexJFJStKtrT76qhoLQ2YZTE
NQdpJrKNgL2MEsosZg6WNg24V6MsGi6hoAQaQv8CTVSAxKYFWpmj/9B+TSfABciU8LCaISW52dOq
4c0ANPc10wYHcBqkbOGiDN93XmCOia/PfKQS/zj/926Bgppv1PspFE840dgmihFi74yLzC4Twgq2
yu/Tm4uSaZ+PoKo3fPw8/lHaFEXidcLs+pJwmjL3qOn4nSuTHHp5y9Qu+UYPdqZsZca8jfHrGrLt
3VlQk4KbsGyd+38cHh3yJspj3i9v00UU92LqWOEFoHeYaSiPTFV+ROQ46QqIH6KaU472pzQTRJ44
uPWBjKhGdlgFyeGp+SUb6rDIhDE/t7bwYTsHVGpRxOrebdlDH2arIke1ebhvewhu555MGjMeGp3m
yE+rMS6fau+UGWhgWbcYAFylv2N8DAjkbMBr4quRx/MIgcldKx5OdduzmO+5864NLRLr0rxk1KFP
zOg6hvO6gEv7HnEsYtIBmR66ntUHl4QWMuxwN2QpaUQfgPsxGqaHT4Tboy0BfxedSBR40rmjtvQV
W/Md/BQBUFAjgWuPWKGAhXaxYDt97tXoJ2ZfQGuPXGSff93M3W8CD6wXyvq9W6YnEh6ay4GoVE4q
0ThhDFKdE/8v9n5K3Eefxz7IHJH6bw735rEfloo0abU+AqGZKyOSpU6Ruw1wUZgO0TEpAEAcnuiM
u5+92dWWcjaD/ol3kR0MRKh5SRNHkpKb5x6qZbKGlsaqCXYnp16zI7ACtV/KSjls7C/wlZrLQs3b
VnvEZiOzw22NJ0+nN4o9aC/Px8wMknKAzb6DDWoiynIhKNHjiW3wj8bu0tqNhhiW/djFO3xSok4/
JdONs3CaR/F6j0NvwcvXV8CZyTBB0gRaht8lmmaeZgVdpxOSmd7rPg7zmTaGX+9/3QhCQzjiSu1S
KqNh+0+kGiCeisKBmjhdPGHNIaqKL1Un2bBHCtC67yJETjl50z/+szFeYX8KuufB/s90+P6r2h08
5C7Bz8vwp+BUf8/2FdTbrvtbMJn3t8uEFHVUQ4g2fxukXUDleAKu8Jw/4tB953lCPwxTCEAA3bgf
AvHMt091HNBkOZ9SOPhJcrwBnEtnhArI/q00dkZXgHnIK3pqd9Sj60mvxvF+wzl7CATCKOkdPSRG
kv5sqdkTMT5mvYZKBOjt91FixX/xTM4xPnRYomf2+iKO66HpNXISIcudUjXG0OqYljzoMmXLp6pM
JpkBVmPXn4k+wXnyU9ewUOedccDacpkQyc0oUk+QL85mQ01NaFB9dGJeExwUAwCrcAzcJzJJMhDS
sVrnNiryoN1VeoJlbHoAXcTI0MOCc+aro1gsfTdh3NBEFdcS1/cCSDG+yvhXnJy3r9vUZZN3lgku
MplIta0CHkomOm8FFYuRAGJxqLB+63M/f7bvku9/3jCORxI8QATvT4BpdhNH5Zcv6eyOpoGoMoZo
wI82J7w3iHnP+eBHlaUpqF2TN5L4LjrFPrXwR2mI2KTo2FOHOQSBcjFuZXG1Uk8H/sEJ1FSRIwIU
pNc45xOM8tGCCqEZDaWTh1UhtO9u182L0SEeW+rlzP4Zw9f6jGCOBbOl2/32JsrPJjJxOEhtMXco
lUXXPO1er1APVr+RU21LTJm5CQjUb/VWH9LBbcw9qzXKhxnShB+9zynv/7vXz+3/KS6q8mIs7q/1
Eg0MikjttYjdSMfCph3mFjJlgWEg/dScCnO7BRM6k6v+XxNfaVL0umvaxWPAPzXd4wHzItOLGse9
s6cyOBtef3zYL2wmHM3IxTauoXb5ox5lk3nI7nWxYmDWtMrT6FbrQnEHtPOvnm0/vxP/oLQ2GQ73
nKcSn9Tu+OmDSvCSSpKuh/1a9/Il67BKeimquTjdxcO8Uwqx+29xDQo9M4Wsr6xPkcD4gFYrL/WA
OFpKHee0VlTnAWkXXNReawV4eAPH55ggeLCjKURpXYNEKJp1XtUZjr867NuhTcsI+xu9meQkQ0WK
t+KDjEhVTlY0M2ETmX2wXtFz7sgR5zqWd5iZBBPd++vbWO/poBYJ0OAiwA5AtvweQKSaBQImSoFQ
fZb6Uf1PCF9sIdwycGkFx4dUAew24ZvBywTsEBZEGsOGz7G3VqlLcj6ZJEGCEoslB0tQWGMmfM8I
0SaiZASfU6wA4SmaXWaUJrIya1lyzOsBFCsk7qF5j3m9Jn4f2NNmCBZ08mw2VuXY8PG72iFyfhSH
hrWKkPE56xAKLmyuRR8nhSefUlWRc3ggn9f6az6mRpSLQBDAEXOyi18yAPXTJakvAu55VvFubFjL
mPy7aDtxcHnFLGO0wYQCY2WCt6e7ZbMw7zEyEgP9N9Q0GCncoRBRyiqxjfzz9ldYDSXctv7msCa/
dTcDOSFK7bhU2TWputK4KpYyDedbFglMnxzwPInjXGJa1Dhv67ifolzyDC/0XC7ivvKtTo/70SUZ
Bw4fVrP4v5xbzhkf1XtVHOqZ/gu3hc4E01EgVoB5WIwq95b5VZI2YZnwWvAkMDb6RDJ0J6ds/h2c
f40WxMFinwrowbeIX/bCdLc5g6YvVlZqRaxyL1xXBF7kuXGbLA9922vv2ditf50MLTYqML/ZboMn
wU+fC4BGNaw1cOj/PRy9qLh7PVVG+XmsKztnNtoSQYmXIi2A4gRJqHYlKtlKsTW1WarlJQDeAWTH
d2UXmOXHsRnVgnchhRvQiFR76HoNb8BZO3amJSpjrHnSDzzuN4FRNv6JPFF/ZMdBYgQBSlMjXNkG
b2TCTyDnwR/4rfNpAdWloYqGWpBWlfAz+fHQleSkW0yfgfHJqW60da5wF/Sq0Sa3vlvUJTnIuUBk
TnK5vt8Lxy/FbRK6/r3KDc4IxL8fl/VKxtLqwlCE6ALlfzL7yWXywFSBeYx0Ly3iKSsBjQsR2FCF
mtW4FbFt716K2iO705iaC4bcojQQ3tEWRw0lYqX8QktU3+63mAWX3b6XqVUsTDBJIqdUYiPslchK
MJ6IOCm7/WOGoElgsTEeWkPDjBjjjTpL4624F9AH/5ueLO3sjpp0lpn34tIKP9DS+uD3FnhQrY7g
K13cmdR5lcFKKkG/b9kktItc0b1UXEPZNjSzgIzDWfVHDXhCC0dbVyjKG+4OUOTF3mWhI2w0mn6s
dU8KIY1aWjdIId5NBOn2jeKgKKt5E6HoHTUNejJx2qusqty68818peDa8Eh2qRI2isbitGgpTJr9
8D6ADfvsxjxfED+fIyjQY9p4XyDEGgtRbO8CC5T3pCaHJ/AdmRRZp4QF1d0ZiFtqzPK/w/35/UZA
A8VdvhJ2ooOTDzHaF/iRjhdHnQusiZVG5lUbWMqg2JpFaQD4z/geua6dLJhwdW6ZyEEnaEUeCtO9
PYA8gNTlt9SJc1nkCI2Y9Q6rFmnk4gHuvl4IcGwRTvtrg2AP+OdbPNHM3DQxhrDYDLTK9fqytKAW
vQGtRCMT4xoA07aTh4AahMIiw54TwhlEBFrwXOTpjb1uhKdP0hzqfPEcr9ZHQr7/Zj1ObOj/Fn+I
ZIHsiylIwlTsFc8HpWE8pYOpnPr4f6Q37ifmZ2tmwtAdiRWphjbmn2j4jhrpiOx4DWRYya44xhjf
PfgUW4Pa+ocieLmECH4OG/zEcRUF4m11E1+kLog5fcmDrcIC1ujFdSg3R49qLIh34rdzLhBacYeg
YiZgqhQMp3G5rcP+K8KKsjoAFa8+5Ka8LfU8OK3I3WQhzhENUcWqybbVyKVKrjFi5wDwkXV5tjYe
RYEowLiqonwVUCSvkSsPU+sRMDx2ytVsGnBobCT9741wWmuR8Xt7YNpNKVBnhzFvqz6vBcNkdWLZ
4NjI+wmKellciVI07rwoFGqyxTsl7Dquy/Usl63ubA1wyOEWz3cA5uSZO4lkLtCnWzr8R5RMk/mU
rn+ejjo//6bPnDOUizrTWzuqAHPw8W5bZhYif07n/lP9DGVHkW/gWxyfUSv20PaC89pqIH6gBr5j
DdTfzkEdV+Cci6+0+hHyuEkwkRfdN4kj0v7SVOySawxAd9fn3jKL4FZRP/CzCPdRMqAQ/mDN+OIG
rDrj/pAKdrHuX1UzCRJvK0VoCdwE8mM/O9/UzSHkM38/rWD8qHG0Ri7gYvRHYSB9VH4evJnd9y21
kzyQqj0aaqFYBirawGme5bf027N98IQWoFnr1OFsvf/UyNLp4SPNWySD4cyzMuMCa/Fg0q4cttyJ
usNiiF8q8TdAhybACGZk4tqsPq9w7BYOkr/TADxEjwZnF07zwwl8yKdOIVh3O8v61i1hafvnzboD
kcfD5jk56T5zBfoklBdv3hs7Cj0ZzV6eal7yOQCoNgV0rumnuLtC5a0Sr1EzR7q6DfZDr3NyfRSN
PVzPGzinfiTeR2N+zW01jOCtUMwfH1kuuOfTb5CVux1+Pw8jz2SQhWVKTq0UqmzDu9dwdRlrTfw3
72jUMv5KH3R1O+LI2CQp+kCnoBIkF2EjW+czAOhY9hFZYR4ijCv2Um5riHxAsJm57sghBP7T08QP
D4UBiUc6LumJfZZ8J0shR++lOM53BUY1qzA7vtXLAO5sC0u7XHukxKvCt/zoYNgdwJmTRYnDjDVS
VgFHKJqgGQoNuXDAHnh80b4UYvBjJx1jPzoCV11sG0rf6GYAR29Kuy49yi2wDYKPfjr2+ZSLbyVC
BRTyxkXE9tu2Z79cdvRc0YclMd/2e/z7FcUXvx1hCEnveImzCnS4QXhhjky1ZS9v0zb1VfwKmm4K
vyG/VYvqArVhOYQoAzXHC73pH2JEWSMx1rOU7c0rucV9R6+xdlUuLnFn6gVds7Kftkf7Iq1fv8JV
l4c9jUGnNjgg1VWaZ0AszWu9LXScxfV4MdgXbZLGRJyE8Z1DjjY3XkLR2tdh9gs8ukP6W4eRESsc
ETozhEqwcxj1QD4qoRLUZVq4990frTpN/oNx2UU/d6GC689POKTCqhsqqHAL3RTWVM3U9G96dGqf
kdkE6cEtL6RWla0cSbniKN0aGM4HOIlRf/uDCSqx4cCUgKQgTkc/OBTzNpHOw5MQAO5TgCFqW5hR
pUsAmx+DQCcy3yYR1CymqLpmtRQt3bwnZ7UuCCT+2+gPQHJmsDd1+4FflP7q4Fg1BtFqJPcqp54F
t21B73DRSUbTFrOb5mrzP3B68Sm41/5394mcQ+00UCLoN2JIMtxkK6GkgN1rc0GsSDex57G4qdcT
grtid0qD/Gsumnp/OlYKpy8UQtS7ngaEgQKytIKs4fRdsDb13Ps/u4Fy5Xtn2KCdbDsNiScUbqba
7JA1dgrCP0ajBRWapbvY0alA1K66rDkdyrtoV4Vsx7+HSpIginvzpEcOYgzTpwDM11wuK4LFs99z
58GxvkU+7DodD1m9S7CZt29IWIKQdTZ49yBhWbVeJDrRn7bjRC8fGhxIthlfwlqHUtGa70IoOXPZ
OJgFd+e7/XMXGMyPwrZ7lzEv4bt7aI0C0tn/+IIrWRnPL8BQsJxTSo4A4Da/kYPmtV/FwtawMOjH
8VU78iQEQ3AFywWtgL6SepyYVywWKS4wb5HQmVi1Z6QGgy4G2G/9AS8EmsC3TJImh368N2mDPiPG
BeiAh35zwTvBJMXz89PrPcRTB8iWStKrwyTMBP4zBNKAp/ptZN5fQCqqcC74oCCogONC8fGDzGUW
1G6fea66w6PqvYz57pKBnqCQm6qTcHrD2g88F6iP3HbiC81+MPXHzGRNcZHAL93Ql03qZ0ig9DWr
SHZg+C/PBKl79Z0sGOgNBO0dpBViZT9Vn0lI5A7pRytXd1gYkf4fXpz2gZE0huQu0L6dDCKpXNK7
8C9+LFUugi2nds3ddpYHIIZiFAsC+M5Y1j05pN3wzMPEt47slXy54+xu7quhsJnMyIbbzw7xI8L5
gGs/6gmlTwbBGTI9W1ZXG1/6wBv7S3TGKqUog9l6gmtJcsgT/5KzburuUpnFv0fpU8sEY22WxoyB
8vhm3oS9jV4hRqNFxG1JOSaUivI3mwCdX8SY/ikpst9k3S9w/jOt8To9naL/gDkDC2Hser8rKT14
HNvCEs0DKvEDenyFR/sKCqyY5JmsRsb/bwQ2niaSQL7C3P61rsnhG/Aq4HYxsLpxko+/TsbIfCej
AFVIfvdufT0DJab9zQhDJhxM1+N0IBykBrcWa/79PsrPIUNg1xkq40pBQIVDy0UIx4PB5gTDP/lf
2Ac3Ld8/6aCCEMM6VEYg0HBFYEtHurQbEebRdNUe1hbfqYP+B7+ASOwHQuYfahrr9qcnhKqoboe1
cpmUBW5Q5kRFhWi64VwrtFDr0y4EE5BNlEG+U+B9idcw8btTYYjsI5OW6IyPg1yt9gQQVROJGBeF
qPtGWq+oCYJHWnpkp7qPhUzKJFCbYjEmlgiJbuJAPwLuevdJMw89vFTEvc21Qs8fxghaztWlOEvf
GBdhN1elzNR22s0ulxBWGB1ggVz+Rdn5b6GCD1VafPHuVM7MdYVovAKK/02Ae7rRWwUQBp3G6ygp
xvRJgP2cn20UQEXSe4kz+hmV8G1mbdYNMrUSYKaLpSpzui38UHJxDePjqC0KYq/INIJM1o/gY/be
JSnYPaSd0qTdhd9Kd0Y8uOtZoSL2xmC3KCb5KLC8EYktaVnVSyVAEnEwwt2G0Dkf5D7429QvNLL6
KX9+IfkKqkVNOI2pgjgrC5d7O6TLBFGRS2ucSjj3X1JeQGCs6Vo0bcRZ/O+2dPyeR5QvRAMzLqeI
3rkuqh/TpccguVhZ5x+fWOQTMT90KGrP+IxASDKBJoG7HrIr4sFtjRvE/xGaMd2Ge2+Xmv4Swy4O
YGBU57E5gsK8b8yYjfMrpcF2P8Sj36iR1YFrLrttivtgB54iFbAAG6xRle4jvXc+EfLhljRZaMyB
mcGeAxEBw5GKpAynfVFQ/x3ohmL5q6w+pN3akc1JbW6L2STrrv2HZjcFsW2x/a3HGAT7Iq0mbKM+
u5VJIoLISMU/2HtoeWjfLkkDFHqWhU0UaZxMncK2IUYgtBEijktE9Ye4AIk8q+0Qg7i1CsH5VMYD
YeSSXqJr//SmfRE78S/pjkAVxa9/jUgflcGrzjk1HXJREYKGQijYGooyWPHXS8pG0/pKKRRCqrDl
h2sQsVyyCQVSbULS/qHRj4ZzHhJ7pRiLUvYJ5Ulvx0zo/QM48WzlcpX8xMOFxtx+iRELxb4+NFg6
csAlwG3OmQXI9uxhaGRXMgWGug1LcyOqwVd4EZGr1mfeoTHRtHhGycjOpJS2WRH2WLf52DNma8ww
flC+NAn4SFkscBdblne4rsi2FZ7jQQ2oxNZ6fOxo8tEBlqLHUmmmJgEtayM6OVjj09Z3lutEgV4v
w5cMvKMf5+Dz3pSWgrIgXPK7JaP1jIdAnW/h03CL1UOI79ksIoL6L2ZWVZ8f9bKal9H/FHxpdclu
X1hWa/8h8YuhCBGHrxtAEXbbjUDq9fYCV5fuljqLzYHoV55SjdCehoJWzy/tr7LOpuAK5XKKq4uC
OGTU0rqnB1Hbwfvep63dOlJBXYkOJ4jUxRv3iZYYnjhsriAoQEsJATblQuPgyEBQHG0OqfqZU4Pg
UPtXryzjqRrTY5+WqUXpcbcfALxILM0hrmPhxTXnrTHI5ISCRQhu+uxiuFEmlDJ1kQudXNCdZeCF
pDQlsYGy6GCpZrT3rVoTRiG+bxg3rsxqtbZnGn7TTiumZydqoW2klUsl9P/XIk1vuGAWinkhyT01
97h6whzq4DxqirzaWBY0UdMvdehNy8eIYjewamZ4YXV66Ies8wkhUXQhWBbN91Z77Cc9In8eUTJv
C6LRbwCBhJji00+Em9gyh1BYI5b530HSfuiWMpyLyazlwKbPO9P7hnfpJZuTLNMu5kroIHW1xc3p
yNNKvJybQL0z+zQgjiAMN4OUufOR/6b1sGM9vwgoUMZCXD0vEL4mqsvbMPioXqXboHnS64ICfAB6
FCFI0/XdFaW2RrmgV3zrlIryRJCLxQ/ba+MXajglPmyDxHejKyWx6zvHC7TmZScrlncTDIRDOAPZ
IBJM/E/UnaSo/ja2aaGLXCCkACrVuAO+MukNb4+syEEJs52CM7/YMKy92WUpBrUaWV84MiqQSCFx
LSoUHLSvOQ2LLkk5Q8ozZjzdJAGq3vTGQHORbFBSCndgELL3gKjrt3f/CwBznKcQKDGZAJwVgHAX
u43dnx769OL1odP14OyONCrJVjG54E/CjGmYuqcmRvYJiCiOFCcjnoi0fMXV0VLlZBrPddVh7i4x
04B03nzja2muUfInGJ4gI/VRzW64pthiy85cDyQsl5oFj1j9ywHvhgXg54cIMunKXtYXaj9+cPVG
n7e02nRIzrOPcAFSgtW22TQf6qrEtXWosVG/zKdomLuPn2kiioW/uoVZiZVTmbT+F8KWtREatKHD
Mbn36goe0fmMagilHWSzEUY0ewXhR385aEPwCLcaQ0/9H5gAMOyX64GbOPpSTHbZm3aIlzT3sKhL
zBTpURnbPPcOMaXGeIzYIsB5qqwsMn9W3Tcs8+INj0FbR1SrqTSrTlGPVYhqP1rPYaeY2nc53KS0
XNqsZ/uNZSTn58C8SimLsmZ7fLanG3QTA5VhbZXWL0dJsIELkTJVNQm1tsnp97mIR8jvqp2O5Stg
fqpD6/7RllkcL73v2TsVX0EaBLN3WZPKvrsKzLAnib2zAFE4g3npyA6/pZfH2TQ/h2gFQYg9WeDn
Znsn1TUWnyZ90VdUqzhPxS2nubH0RIS+dIfvNNkbDoBIPog7g21nJpoSerRmNlziWOx2sdBNFMEk
07PeFF3a2cpQjkVfXkTICBXX/iun+cD0/sl9vhHdQVr69bUDxt435okGdRraUUV3zHwO8TV37/in
CZ6d/M1Xdm82kFZbVKd4Vt7R75ANcj6mgSDoWXr4PDKDSWDngMnJLawn8pcHyCjC4LnQDF/fq6ZX
ja7ZmmUBZZSPj/aKUr3WEfDiIsVeQLb7z57N2mJs06lqrNoHpFS1W6LgYF5UW0Ouh9+QN0/0HeHg
DUK/l2dsmkpamz0Y1ev7PS5TRJfdVqGU2+xot89Yp9NtqgfUDhxTyHN9/kbaEWgkGyxRwbUFAEPj
DNZ4T5Sbve74srAfz/rebWabPsHAs3jH7pzJ2vSsu0z9gik86jUnWtt1CQj9Nm2x38ENSAFIFrj/
DSYOzhnV+UPsAr+oATk728UUPTicvy5RuxWJ61qhjfLrXoB5qeTEBm8rRRp20A4rKgtlDyoV8WZw
Q78jZFNyQ2B/YP78PejM4OxFjQlpjvFmbXoqfeYWritfn0wLLYca2SxK2DqGXXX+CqJAQFkCr5rA
8TcQDYbuuRjg/OT0nnzU2G3kjLPYmrQlcIT5i6SKeg2/cxMLnLTjMmUW6XDD6TbJAky2AaLzTwB2
eox2kp6UKP4G1JPDufZ4Ap5pOgPa3HRss9PVcRd1+BKJbkpvWoqiHZFo2FfdoQwo50mqrcaTxZqb
1IfDPZRkzES9LcMTrel+61nBUQzMb4yKDAwCYFRPs0bi3XF9iMvcHN4lLzkTNALJv7XMj6JpN/H5
DaalaToP9RwlUF7cXJ4dg8AwQas82jCgooExUPuki236WtFuUQqJkIy5WZNTfsqzWZ4F+sJ8PjwA
scEFDKKH/AAccru6T7qEnatapKNdyVTJr9kUwIDTGd1jbYj/WBGJnOwJjj8SOHHLbmIqE8W7K/Ta
B4uQoIgGklNQSNT5oMf1vKaM4acPgpASPHrsgkXerKPlZoYyjDQgg0cZhT3rV6qtLic2YZHPUdk1
sXAa8asz+nByUdZEX9CsqMNeEecSc84+cPar6rsC6W4ifqWlECBWLvMH+9Dijqrir5Fl+jZZkefj
GJi/ikb2BZcx/wMmr+CNvN+uBXMlynKzq8cW7QieLdBHau3mAZMMAsvA5K8E1sxtAuKxVODcLkWa
/ua/RUJ1rObJJhmhtNZUAd42/xuVXMeY+8l2w3XVwRr60q+ko1CkJd93WVwu01by2R4wDOEeRjNl
CHHcuOF/9z+yQ1hfkSiMcnAqPvkHn9pR9SB8RGGi6coqpayQxDQ/aKe7xMvnqTUxJXw38zWF1W0r
SVU7g5mc+ePxoyBDMYMaqgfnvbYFdXzKMI8wx16JAaOxAGlLr/DCaOB2ZLpHodbu2rJi3g4bLyXd
jSWKqtIWf0CpconDsQyvFp4j+S5UznCCrqeg2/jrdntz7YLChxa6QTz+Rg/Md+JpaXYpufNBvwXn
OnV1ncHnC1T65SDGe5Ry1J6vIr22lOOnUo7a6giPF7BibmpUEn07r41ZsFrEFwFFIsqMnoNZi4u6
bvPPDtwsE0SqYCT40D83V5sqBBYVzgxlDLmU3wXjnX0TBgqamVhKkTbHDHXiKEwgQvhLU+ErrpXi
2eoBMY7MWAn752DBHb/tO6ldkdaniCV2hvpDgp+rY1Lf0Mp/1kw5+tGqWTovVcB3cUk0vXfvfksE
iXQ3HgzdqYOqx0vu6655sgOyKfjtEUuNgMHKsMv8aC7WKKmZnbw6Koa/5gNy4RGoPlaTCVtBFNYi
9FQHst6MJKngCxg82uz+3Uuwu/Tx6MQSXEnYQJLO9NcIZGqvurxktJXCeHKdYVSqnUtOs5wwhdQK
U3bEH5E78ycHycw/cLL9O/4k0sj2XuCUZrMSgDAkKGHrAhsbL3xWOFJKOKMVEepZdKzP+2Pdt6sJ
4D4PNqBYpi9FawM2+HgwacWSiRMm1B8QhjBjc7rPUbGT9YteakloE38I80mELVC8MxS1cIVOQHCx
/oKCVA2Ce1ifKK5T9B4eZsWpSCSIJp22QyBCOY3fYd49HPNQ5BOE/zzg50Oje073STffF+X9J1dr
eSgIfjFf7s4VXioj5eB2BaR1xUl6NtRClqtHzCUnWYvtrMf+iWtaKYHsob0yXeScmyMzkVLuBm62
9+pI8jvIBKbpaWMmhyF6iribgeUskwOVFFaRP/V9izk4pcwDooc5OjKcsvP5s5lYggqkkgdHiC4Y
pmI4QfmUI75wOTHB2+uoXUh5DGeQJ02CYMZBm6oYD0veO68wyzUFWEMR2eRynMNjgRcuoKWPGX2W
93zE5l52REDHXVGC3TtxxDd/wnlAIaBhUrOBJB4KSqUzVIcy7ycW5Kjin33/5z8GZofrUb1Ncw1p
gM88Gt34jZo/fefhObEzyDN5y8ZDWP0JNGPk+u6Tj4kE+G+XktXlKpjdqmz9yBw5lii6DQZ5x3pN
sV000G5E00tv095zw51kX54O0R8Cibf/92urLVu8HbrW3G2JPNjc/ujxuxyi2EmdO0+CFAr8T95U
yfXLW2ZQfgdyzzswAZOA0NMOE7GYyTjVbvdUbeefYMXClva091l7pPkXkg3PMJIgLCRJNlqO4ARR
qNTYt2khFOeltC0dXDTWiNF0dvmh7FaCaTsQDLgKyF9J3fXJidK6bZYypFvYRIx9PrTLQ20nTBIC
mVC/5UKcqEUTuMWW0t/p7vemhTvA4CN0sGpsXdV6gdn8TT9ORkA3wr7UhsmZ8PxZEol1+SdBhjSX
6AUELZpVL3ao+7lGiS6OCrsnPz0B0SVxxpVOI+QRB4SlnuXdopyLK1NrqoE3QKD6/d+SE6MVWYvq
VG/SPpGVgSYvy57K3ZL48s+LQ4pg67UxxUFOOcY8cE5O/rY54UGJAeI5LiYhfP1oColSuW+8sWiP
vKnaZdHU0PAmyf4somlc9xUC0go7KFfz5c3+u9ntJbKIWrKIPGWi1EKp7iec9afbxP7yc79ZlT3p
LelsguK2qvnbPOIqYNpiU8CNOKG+q59wBu7Wj4H2kFROTwBbzvkW8b8ii+bnghAs9+L3JbaQI3qd
QvBFua+8CAh56BPYKd1gPkttLeMXzmuHgxgYlDGGamH3Pp3A9Zp6dbZB9tpIv21fivnvl5Pjy24o
1tzT38OSP1GpPG3oFZhXSckzRSoGwc/h4Xjb9dTao/NNg7OdaTwMgrOk8XZDBJP0n8CH5uBZh7ky
CvihXvyJCfm5DAN2Ubo72+wU8U236CkmQ0SDg6mGlPZai6gDYWuF4BwzcN4L7jDs5zXmBMmZUf08
ZzN56ZNmJZwvCX5uECkFcrTapwPILoIbo1vJJLltzNCkJPPkRm7HM3PxfSlTC0mFR7bNa9eOGx3A
RnlpDKa6I2gjYAh5h/WpzHDKW/Se9HecrCu2DWXZi3t03mCcdRtCQGDWCZP8uKA9/La398FZOcYl
+JtCylzkYstbsbk86/RxVgJmKWOa/WhitlxlBFFoy6eLVwn+s+k0TzqUkYFyRg90k5K+i5nOSvaF
4rDTc3IToRRfGCT2lUGWaLpLhu9Nnig+Ctxvr5QtlAmpFjN+YLv3NONKqYjHQhMu96eGHxfPB6n6
QGR8175V5BNFpYAmLAsvkiWDjUtF5eN5F5PgzIc3cbXIbEGtVoatxcseAwzsONDTqJWdZxBbYgBc
2JhX1r6qQ8W57kmW+ISkgC1g9DtFKCtSQb1+qi/ULrlX94b5WI6gvwR8w/Nu2dZ5bNLZbtkVBuhK
3rV8IfIdUx4YtuPd54YigsXeuE1nmZGGxol6LQyJRca57jdnJHR5/Akyk2X+X7h4Jhc9VUCSZiTu
xtuK6hZstYAT2dxhSnCQZ9weJr2xEt3rKjgmvFBX0bIBVA/CNURNoU2vDQfSQYs38RrEDtuSqYsr
Ko1xHHpCUK5lBx8j/4yzvLJ9I9ZaR9s84IKLbl/nfIEsYXLvkmjQEDu1ifFJ01Ikx3VP+2IgDDTd
2EfpodfbYnJWOK+nEEmD1WdnVC2CXLnjHG1YNx9xg/5cmI9wXJ+TLZnYZ6+CtZSkh84am/z+uYSx
X9vRqn1h/g5XCR1engK6GTdFm6Babgktgy4GCZmV50r67EObfBGYkFMzP/n+a5G+EJzDfDWhx2bg
0jUK5PtkzKy+DH3OuYwdOZB/Nz+hKwkHtrsD7bPfOesMHNrXKmFGUy1Y/EY9wO8RHbjXITVDty/Z
mbz0VTQ0IjBr/U4VUhm/8vIvnvlrR55lrb+z8Cz+/qw4PNVq3TH4vVOslcAh5qeLcLKqQ3g1B5/N
ZnKCMyNDezfhI7Wcm2g8i8hsK6jSCzeeWilZFTIJeq9EFcqQ+DRjcpnwu/9jYSDMY5kG/dII34WG
KPNExj6g58ajwj3Off7rokqKX0HJoqlBuKj/9QUz1qLB24pMvSMcxtAdpep4i3KWqt4NWTcGeKFE
h9Ge8X9W9VMAqWhgNrpuCpp1Gx1SZSwoTpdCnu55e+PABhN3Vtx+xnw+tT5AcNJyyAE75I269N3I
OT0gsHUwDGudfBNKW0i8OPbajH+fXTM9hhPWUkdm0vG/3Yo0jAqwOP64bMmzYSFjUAeL8/W94X4z
UO++8kRo++bL/QPDczHKJZmNcGHY3SMvgHBRXJsy8kOI3uW/6HdrdLQso3xz8TIAT0jFzUl3u4JM
3lKVfSryBD6WyIMRPd5ANWVVRXEkDTJrTH+l7k9F+pvlsDuWirDv9/KS6PmSkSNbI8PkOBZFCbLO
CWhKrr2x3AxHOVymu5BstNRyS/Vsp1My9ebJcpLV9XWh1gWbBW2+6PKIl+rYz1OsLy0ueLsJrLml
OmICZ1cZzSAhyIom3QJv9nxMMvOckebgFh//sh4El1rimr4dMubECRBKGsMbeoJcN/OVr4ztKw+2
f9bq4fA9wXVVC9R/1RfIV6KgfpXYH59xToDmplKV2Gcp6QbyJj0+1PQXveZzH7SyTEEGvtStJwvU
IKoSHJ9KGMccpS8n9eaa0QgcM+zpXuCIxs7MqbH1gK1D/aqSSdPFefofuuMkFeGIXS6O/40ltkDf
26li/I3S1iDutw+Gsc+ejO0e4LhQ3H5bJsz19bVNa3eDuhO9DUGkXdg4yK1moEvQTDUlomtGPQUT
LCrzwGQelISKFLW97pZsuvOIg2b1z9YD2MAraJfy+99FUPB4/stAIHfbz/wstP7uVwF47ImFfzjk
ZFykROyZCUvs0h2+em0sPwbiwNLYcdXfHdBgJnM8BWX1mDbVtacq4HWmTDlAb0qsDqZQNOh3RX2c
bZT4/zLCH1tfXRdh2KRvMZmX4tVYh5qk3PbKV8CyhI0BxKnSQCeytt785M0VW8AiXDVBZiu+wHhh
/1jacz36AvhYqbUvA/I4lIggEN9ALD9HSRBSnhvjEObYQJqHcAK+NJAmn0I8sV2zIE5ygVWDFs7A
/H+H+2rqLplvLfUUdsJ9Rj210KCm8rypXoWYM5fn09LnGp4UK//rD9tjW7MHRB5RnJZvtq0cTlXu
2nnmzdXsQ/3CX1I0+tWf6/MGlDMAm92wJB80HuSNwVJpyHbKfHDMmpLoJPXmDMKoa4nF2dm/XJtX
ZUUDy5D2MB1DK2xnoqO2XJ7O+5X/szQBDFLVRyKcviAA2UbRoeQQwzDZG+iGhuPX025kgLIwLG1r
fSuqWFymmGhuMWKnU4oz+HaeKUb3XmSsjcVriHfTkcpNCC4UDof0lmMwvtMyiHemlMztvFUhQJ8l
dQEWdsuCVvUuEaq7J1VIHqcxm0DVz3bWLU6sWR9elPQj35ZTHcgx8C5d5OOzhk02+K/X4Ia0H1xl
NlS+fIG6gaHkFWCVZkUK0VcWnohs2mheEiGITvXkF+UtXqbCJY9Nsaj24C1sBL7MCTvZrGWCixIP
bzW4eO8D701bpEVSKeruI1Lgn7q7yTxhC7z/k6LTZH0E+xsTW/mEG4IRxP61yEQaUEvLJ9hJGriF
y9OxmYrOQ4fJdt7Bo/YO8IMwKQNDAyQTiTvsY9K3THXGwj8Usq8cRbtHsuGxIV/5WK+XHxhWE5WF
z5uZ+Td/KOu9tpYGYXuSkhk2tVpLTFU/S9HqemCe4xqRlBhqLlKoBnlzoAenxBJwbewcs95MAMFo
SvPO6sGDZt+V+VJKzcA5VJbW/997pB/zkCiE9uhPTJ4MU4jYKKtFAFlJ/AOQwVdSmdOUT3bFgriY
bq6Q7RE6Tl8kBruwfaJTvZjFOC/MFBqT8I7A5YYdZke6dexhZuO2O+w2ifa/hRcminOu1vFsj9z4
BClVYN+P391m8bu/lXeueuFBoZ4b5qy8ZASi6TIIu+o7wQhiHvFlFtViIOBKZcYFuL30HnnVeyWR
DwIY6QxO2U8CifBkoANmuXW1ggcmRmAM+zq4EMKOWFz7ab5H2Ryk5za3UjwQTCdi9NDXI8/YbtBy
QxAMOsLbpIDFBFwKiEYVW3Z8EltslVOFV9obSjwb8uaGsuwfEPlxUE3DWEE4LWVHcJJdjQsyed0K
8+5XylsQ9aKj78wopIx8vFJFvaYRdkZBfFmtlNQ2cDNw6gbm8ZOreKyWmY+31AIKhkyrnz6ruXxS
XTO/h+bsEUeJ4fOXSauqgnWvXPm3gyykNMDPYDgyt+SydD4dkh4vdEnl3DErRfA73OfUlaBr4aIs
3pqmFhi+8ayfsFgYXo4KMn5MDwAAkPh1K66N+ajWfgcvT85QrIfnunddaed96Ti9Aeqnbo8I7wKN
t/A5FlAcwlzD5ONch9ruFlz5AxtLXXmSh6O1H5gx7U9HxzghxD9J5hFuyvDImBGr5ppOvP3EW4C+
8+nPlNuky7YwX/LEAzmOKZYjsH6oDA4UOkBswXb/QGhjOcL7TU/idQ777ishDxj/T0yedhl8xHqD
mgm10pH7sDIYA3crEax3Tyz0R1QDlqb+q+N8y2n2lILrIOzYWDcLn3mxDY4c0yXhHxxAe0AjhDwO
rYy/G60e5sp3YBpegY3yiqwbqh207Aq2zzcDpr3PTXjTmcO99jfDkhgEHuOUAdRdQItaDtlKQN7/
fZjqZtXT0Q+BqQ7UGfK8cwPSfFN73gT+r1csMRmNS66meuiDg/uEGONJPAZhSOpmxXTjep8IZ9/s
OaGFv49paux2AgTFhNhtlDiRN3TnQuIiIhPD/EgAYJfhO+uQc6t7lVgbIb/9mIJKhaQdW59WmgVP
lRilxrOfYlj/+7Txcyw+5NaD0gzBu8HLQ4SR5u1ZrI1/Yaa1QZxqBmkLaevSnP+rDC0846InxVc2
5LGURsHg+t0RxNAHJE1Y6mZs7Gk3D50a9G8XWkyltBIGBfHupsDS9OvPjo/qXUVlHoZUrEiMQwms
NU3ttpgWsUMY24GQX+vYgmlmTUH6kr2iJyN6R7+VLvWCovt6XnSQcBTSrndnhlHbn+HfXwBitH5X
aibDlWermEtlwryHTQe3HMAlU5t4/RY7Drcgg12JPvZ//loQAQH/lhDviu40ZSx0g7W7rJ8KSqzW
hdzZ0bEXW39wKB1qQwlS+wARVB5s73BdYsEfz15uVfGY7roOe9nuvipGZ99Pn1XgM008tnE0mxAk
s7VMODCMx0G1p5LmSt6MJVkXMgqs7Ev8HCiNIZ+el0EPCchEBV9/TxoZ68KdbG5MgKim7cM3SZhx
3HNAuFPqxUX4Op7PQWZg0uGU7A6ls6/Npq1uE9/LRFmH+RuF61Bvaw/VYCuQzKWqWFnVMQ5TiOvB
vMxiglc2FkkG2UNr4kqC+Q2xnN4QLyykgBtO+QJAJEjiD5DwA1qwkIwkIsQyyauQg5o0JOdT7Fu/
tcRWlUBt2Wk+/eFW08Dd6jOq9mA4FlSS4upTmIXZn/SMzdysQU1JUU4DCHemrsa3UKqpe3mXMTVg
FDfNOHrEVgqTGunn61hC0XXaHoSvfaybILjJvMP7CWdh6hAAU0AvHFKGPf/KvhSIUvpx5mfCR4Qw
WpyCz/UVBU5AZawMF5ARDoHFt9ggQbLls1Jw/AGYkXt1C5jjkxTaMx5KxIMH10G/AcZ9PEksy3iG
9lZjYl/quLm2Bp378CIVXNPMII/Mi/Q+11VxkFBB/Iwu9E2EfTmUJfLsvzR8KwrryaAnZVKW/dob
aKdRcuNvDgP2iOzJBsbTkLDnLD7Ml+6qViERISFdv+4ZlZQSmELDpQXps3ZCJiMDCOoldNwWn2JD
IDX0707B3/xe9fwkfsEAS9SWjGIoV2j1gjrCH+YVf6+Hk/GqgYub9PyUstV3/Hz84Qdldl7w+1tJ
2WKkoPmXXtsEKZKV/ZgvFigrEXNdbW9DkVJxfaYF14GeqB7Jk9nyFvwNHbK2HggBRPma4dAK7LU7
eHkyGVFcYfFkekv57CoLPHX5WfDRmgimVjD2zYMsL1Djh8fi6vG+hRA2FI81v1pGgqyj+nRDfBPN
enPbi4zdd+ArvdfkROU2xHLz933E5T9dNrjBnX7z325j79qZaouPleAD4q83Q5CR+zdf0Yitk0Uk
4zEe7iFdtPM7Db3XboLY+WkV3m1XR1geSy6+wAGk+Fop9lrfOfEu/aFTUzM1/Eo6U7t20MxW06T1
ejgphf7byeU04jAyhYx4KH0i0/NdFtazxR5l2UWe7JMY44zVtQClG+X9CF3vn3QPz+vxwIMhderG
/61+sRGtX/s5RPyzpQV78Ra49H+hiIGFoqgsykCx4b20E0/u6JFnhfhnkQScUP4bPybrdrFn5eYn
v2qBSzqqxJLo/WjpLeDOteBl9oCtA++6NVMOeKaa+2l2CYaS3cheKn6JslIrEy+vnbtrCD+vXVN1
twyse+3YG1G7np0PY4tYgedCH7I04lBIJqz/4qXOKm0rIzKOdVnJ4txx7j8GIpVsJRi5R1tuiYuF
bXg/M3fmM1fs1WZAp0V3Y8V4rknF+Gp5jOL5aMa1LLR+SrSSR0zmkWoIg6EMteLdbnHxSjq4PRsF
U4H6wxGM6lDh7LYXnxOr3M0DVnmtIr0Xl6D0wDy/v8rqLKP6X/vqdW0Ll8zmeVKTPGRpBHpXgbiQ
gD1g6zycAMVTbkXm7ST47dfvDK+HoEJy7gvdCKpExH/rkuC2aRtW5m1LJRCRParqIuzmEvUNJhqc
/ji0Z+tqPzjW0iYsyRETNlKbHP5whoNDFTVsVuDhxKJLJ+G5PHtXIz76nXd9uw+1JUAgogpDVwgx
GW9Zoc9FO8b/Xarpvgg5ug8l9o+lBh8SOt1h4BMJBWZU8lD49Y+X9aX5uJoqztqmf7QRo5ONV9BS
lfGcvRjQ5U+e0RB9kavEeTEVCJfzo30mmKnvzDogSewJpjilNkKqEwhVeUK9RQVS/jQuwwz9v5RK
iQ45AFXxLLWLte2OdSpDytCFPxh3xozMHqQgSi9HZh9tMfvbjtkCQDeShGAWW3Urgx/Dz7wafHbe
RMhVxkFJBbLMEEOdUGijVLmJcg9S33dEo1HlpE2BWno7ZMMgPKBP7ufjsWEf0mLgkGYYlNJfbgFa
qNo4KauoYGOZGzLF99SN78QqxkzlbB0TcMhjLCkXPOrlBbCwKzwYKEllrJNRoqTLvRkHclWUxjwT
y0faRG94Gkz14/AQ8idke1YDTHmSaQi23Bqhn8fXGjKnfZpGmjdI/qm1QmuBtg0/7/Ui6pe1qYIF
axSsJ+ubRvqKtfPeIn4BP+PsHrQfJrWhJcQqcUEckVarUesTbfQ6ENpFj4CWW8ZzSl9EReGeRXUa
XS5Hf11nl8B48DdQVWXmENgmazfYpgpSEQaVrUVZeThKicrbWPRA3WnNY0reD8UwHYfxPeJBjGhj
+teOBnihcNP90YvV2lAkDgxwz5nmNwku5NDS3x1zUrq9oP+Bfq/sh/0Z3h9+BqYzhL3cElltGIn/
Ntj6YH6QSSGQXYTuObdd4aNdFOCBzYhGKjyp7aF02iJVnWR/MmgCeblLNIXk+rDUymRkr2pBUdqd
h8YZUnJI74Y4YLbnPTWZtZzJ22lAUM72Sf5lWRI0N1tlJUALgIogQlZj+AwVGut0XoiNg+SL2ITs
Hj7z/4G0+cMHhrQSVjVcCxTxpDGLTKHhBZm0nPTwqN6I0gNFGDQ1KiMr6bnstcnj4ns5enkrn78y
i6VAbRQJ/DeZp4iFrKbHOBctM4I8AuYF8oW096fPt1RyU1fFL+uhG5u93U2LSsKR7uWmqgVRWTRP
GU9frhDnxyjsoo2eZmUtBQRXLqHFpg+uuz56fJud3oWJ6khQeF0rTppy9I+Yrg50ZwlfhPA1dhjC
bdeytxGJqv7SqAB6PwJVQKJplVBbBU2YLf9cfUzoAZN/Cm3sJuz+i99+OaEwcek3xS+suzIIOG4N
+eJK6d+Bm38O/Luipw7RTBCqRUI1wsxuRScXqFPYqqi4TsQi2xhoTUoh5SYb6gzqEOV1aOQTgYeI
7rv1gsGCiS5QYwR2ZdoW5m71cIw5zeBNFHk+HHXxsYaOhF2ETQLc4oy2OoULjakk8IHeRxI1IvM/
UT2eWAgmlkomDc1VkWTSYbScTQvVUyIJrmtd18K+UdneSh4hVicIVODA6/JeUa240yW6eqnEevkQ
u1tyY74AhFNjwnIEtynXYcyXn1huegSsgiG8t3pK9uSim3bDM6OT7wtNUVIjWyJs6egB4Ne8cB7c
GM0LgOpaVCkAy0CeLNf+7hLJDySkDBHxQ+od7NnvTEJgLbrf+qRraKJSZFibuVR/xkTdYgblJkIH
wdUMCpRY+72rn1uz85n2EWKrHuNp3C2Pmx/YpWakCqPsVCGiNGF9w/Ynlw4yPMrU3TQFSaZd1v/Q
prqU4RZiI5jtWrFUsK9qeA8zkd4UFrNgpCBCnzobdlkn9vI78sct2pxQgV+ND2ccoe2GaMM6mg4H
GNS6EgbzZue8qZBnZUfb5VOKYgck6TUA608eCss5HOe4EX5MTk5mylH/9UvLtKI2709CG37IQt03
8amo5k/HbFfZNahsnA97JhJms03vxv7O09ryV8gTOwMNR0+CDvyueKfZTnimHpkwi+dQ/vAqM7rx
bFE/lQypcWcVscAS6Gs9TSYPZB52Z8N/72bU+i92gx48SmK8e3N7HV7GTiRtMbL7GvQ1iZMz5jUL
C7oEJYBgN05jPoZhbhZkdPdz89Hxt/PE1M0YBa65vLesUZVGe0JZRK/Axlx/dDOfG+7vMGxpMsvJ
1JLuXWOAxNAWHWJC4D6LYrabPZrAkCvBo5+qCyv3tXsJkWloj55ZkS8lc9Nj5qswMYF4pFdW9NCn
FfrrRIjrYJN/RMB5U96uejVMaSKuG/HNiwRzmzQAskldCqgLp8s/0EDSsmGh0fYf+ZKetelfVy0i
TPVF5XDb2+dzA+MzuwJocri5Sl3axo7K4HMkV33ZtviOjPa/0Hjz0p4KyLUfrl3HkfbazS84ul9l
dYd3vVojYVOtt65fZU+m0hhwVEDB2VI58ibW/qZH2H3nnuweEU6uzG8FBT++yXoj5dsyGyvSqXQ1
hM2Kb8+q8eSuqSeEJLizaGE6mg66TZOrRDw51xaCz2cgBTbK/hQmtXGiF0al/PxZvWFjLm+HaZ2Y
rC8DD8qPg5bonKVFNyshYU7p5U5039P8HJsa5kljF4XQGSUWwVMrYWzYBUDWWyFntaOVy9kkU//m
kHaBXstycKZKXoaKuHT7mLsrxhi+cCK+yzNQ2mVTXypCZmEJy2a+qlb+iwmhP0sfsz34UDSjf8GU
Fo3G25sFp9wP7OyDVJwBPqDN7lPWiNrSN1i8Ueg3IlP1JMhefizfn8iO9357XIo2c1ZCr5AK91GY
YTlKXM6WJttnlNdQUjubYuKnwvdww7siqGWj6jNp4JGXBUU9PwxYVwsZRMdOqzAhAPk7xwaXjHWa
6vvhcUXvpYgTbwV1IiZziJQF1SmdG9Sr3agt8FXrhfguHvAbN2aPybW2jRI7RfK2ArWWHusTxyKk
iojabTJYObbf02dAIzkKlM8PYIsI4sA0tbnNgtHgWzxGC5+RYocRm1YtOpmr4XsTAv4PyqyqyRM9
c63OCZqr+BbgWS9vOj2dpvege4fqN8hUwLGkJnSgFMjteKsda6yVCEb+rngoZBbiAr16kznte9bV
tFbreRsIqcr81xbSTDt1DkEE/VeVfi5305EQbFmkVCz06s4U+VXFewzqFiHKIpDbkAMcdYXc9PzP
1tkINv+0BaEcUuaZy5X+Go7VfH7D72Y4BuP5IUcLGYLSw+lauqX2SScdPO5ZF8Jz4wF33d+RyRse
WN21ncdVgbwVlD5JBQrdXoFnpWtZFF8qxC7BnBnrs3aifFXGcjyaZdBpJXP5erbp+rz0HxFlF5KB
hlIXoOF8cTNhKpbz7rlkPKEYUjD3fA47aAC6n8TEqjYjgROIifTQwZwGeI25kg/GlZarPSOMoF8O
BTfTAUdhgeAX1DtywE/fq7ofxpGr9rKiqx5P7SYv6ril3rnMlIgPa7tV/OoCWr2SHAGm4yXCh8we
1PgroPvclxWjDk5N0mccLEVWLSLzEvLDTfNQ4KFiPVZkbdNCuupPk1rRg4QSNZQNxVx/6A2xZIah
j3z+K3nmcyFnkIIYFIhFbSQbYXmf9BVI2w7AzLUUpsVbc8vevp+GlxAwjvH/aZ2CtdyINuRBpxi/
pVyLaPMgPoxKADoZNsqEJQB9/SaSNkThn4bYhckjgFQ5DNrjMh78BQT9DGJ6kkKMnvoHOXp41JGk
eZ3E86jy/PtJ/hOilM1g2yPMeos0o/uIXct/ZvsYeQAPwvfWKz2fzfyiue1I9AaIrBgpH0izcrSW
DCx6MaH3KE7OD/zo949GKw1Iz/S3HzKXTLFJ3vpc+ZzSUCBqTYv4agqbDMVhbczzMtY1i2pUzTNm
kHqeKgmUnxZYTrQsEBeNsKUdEuC97nT+QNO1FYKvnUhua38tNY5U2tWfjICHwmPKrLUGVOiHIe8j
oheS3115d7QMT51EqtkQHWAs7oH8kMqHSsdnmfl20omLAbR6lt87qhlPMPJFrIM9aCx+Tiv3/DC8
crUN3oBMC7rmabQDLw48L6ifZxFVlVyQ9r5QMw2ckDHSbZ4nw2u8eQvBuFbxr5ghpxJV6r+oFGLH
vOd8VGuL+dhHT5ebO4Pm2ryb3uAY2z1oBfVAlxWwsA6517LQIEYx8M+re9cTYeWS5kUhAr2TRpsl
fVPNbyULWaMQ5EhOF7nhwnKqMGdcaVUXe4LnVKM03MM5vqPOPrl/i1CGiW5rCDZWpdj49VFSq9GS
jPLB9v0hACKNpiDEd9jmxDo/0rJlHhUnctbPhTCOCmNnTvJAZJAtDdy7xE7UxErUcjl9Sdv13C7+
3Du0LOvy0B1RlgjvvL6NoMNbGfur9ie2r7GdFlqZsIr543dh9kxcQEsswkST09c0uV/OEYd87yrV
Puvck8yyNQBipv6H6wgz9hRdox47DF3+3sCNfhJrxgRLBMCasPd3wknFzYQXzM5Z2Nk7wINpfPrG
YeXVPwWbbXv59IwzhlR+OL0R4sp+uJY9Ttpa0tOz3zW5241s720rKOZkwnffaKCTAQeQ0IAhJwLS
vZ3T86eWra1fCKtUksOqVwgiu9+Xf37hK5xX4ZTluuaTqlQ5bIYwzmDbYNnfTvMR3NbGa9/zHz0H
nooK7gPUKhXxBVPNmGb/tBuzvMRxcZOU0zFVxOy9hZ76VHa6bFyqd3aqzRNufE5eXiUgBK23YHfK
IiVG4Emj6LQ/NrmtBpEPypW6hvXyKBsBmHoJDAQG2kv9oc9cLFgvaaY19JuI8t4m+Rpx1uoeLk5R
pIg/dRCA5bHiWbI8R3y+t59WtoFjr3tbaqKWxc+jKyp0SlvCvdyVNte4duA6evT6r5rMBMzaSrIV
glSRY1iuJdXZMRVGPWE5SglouaHcgfTPc9qI/eb/CVsle67MBM/LrksGZys4WCFvqE6+FZsDiOqC
0fDWpAwfyoIpt2Aa/aJc+G/SKaklSfZLwcVLu9fu9EmTUhWJEZREQOl4uVF8/+A/i/8+U4Y6Yyog
j765faO+/CXzjN2ErCMlynmgQJ3drZjA55fr4gxBOg3O7r86Lv9snd/VF7I/e9KNLXXuAql2OZ3m
Nl1zTOx5rdS1uSV39q38Zmngjx9WX6KkAXkFWNYVFf6cm2w+OzKpECFt1t50eWsy1CXDJ+d0iGbl
7E72LMFNpSeDYYilDVVA2rVEuxCY+4s2+mbtLQBwYQ0lr8O7RHaUC8JXr+pVy6zLy++82GT7IrHI
pmfGAgM+HJw8/eHbbBbSclOSIgMqkswIZDmqLCTLJv3tKy7n77MQqj105o5tZmbkH+PMIiI2hPYD
hzyZ0JDsgzcHCvfU1kC7SHzPplVsLqIMICd8EIfNQKw7mUasiMPhW1c25WyjXSYnkXwlj/4MPpFs
uc3IhFxISNvcBZPDxWWPS0oj+MHjOlxn0OcO6tSBBfp777bO8qoYff7Ki4ngcogFlWh4nN2O6N4C
vVe+V//9lJr3g9INMSrs9SmBni5jnFClc/wg7sQN7e6n9QVI2K2h6Sqyeoy3wfUfdql3fNa0O+/J
L374gQjaXskINm+v7lYEdhEuv9Ss5ywnjOuG2JNtxC0TUhSGpLr8Nwteszt29eo32r/wAoKCAhlL
X4V5ig+q++A3V52Oa3ueOECEqXBdylZgIhTkt4cACeXsS+BbYwGTTji+C1+UHZW7TQr7GQVDC4iq
m97ikJMIG2OazqF4+9GOqrY2ozR9Bt1euc5snDoZMFYLxLePH69LPVtua7ayGK1+mq0nQiQJq+Nm
3bfk714ztYvAKzv/RVlUQX1y/AV9OMDQzWCoN/vkqzsPNYUWHO5v5rTa0hTZYFcIOWYx0CUlBRt9
GboppDanBdlWPIIJJHyeZsF8SfPThxjVLIiUbCvjlg+evFLvPKmI9AWkcDOi3YjNEavy5PbynUPo
zt3lNJgrcMv9irJ0tr99xGY3FSTNV6apbe18d0nRX+hdTmuaPYYR30bLxiBtkT2vlywvxxT/WE8P
FGVbnpdwhyDrrbxwoOE6FkVMf9f94JC21YxHnk+YSVMo4Fhje3vC16trVM1xkcCVBCAGqqvBe6Pk
fWV3whWQWoJWn19B/idv3ejAKoZDEVPhGqHJ2/jQZvaG15GxQnweZtqe4h4UMimJ16KXqH1WoBa1
0kdGaScrfmk3tfhweEhAjB9TdNL7uWLFMnpg/eBvdKMuxd5M0TVFi8DitzJwnuspI13Nx3Hh2Myt
OzrCtMVFgalNWjEveJnVMhh44m5vGcT+9XXEArm7VQlJ1OxQvogw7TSWOaPqMwLG2Lc0G87SNnpQ
WYkKeEkGhmxli7+dCNV2g/DsQfxCQGUCY8+AYo5JLPIIDgRqaY7Ibv40WJK50n2n8Kx1OY+0dTRn
xMqKrU4iXPUMtE4k358Ux6PMjnzgcUUjbENdqeI8IfNEb4oucTqKxIdS3QZBXxxvwVOgdkLbWE8n
jC7nP24W0CJyVhlfNoLaCwS3E5d/V6WjO0SAZGDq8o4kGG/5EqH/amCQb61e+D83/MPg5P9xubls
67z/3FbG3AlNgudD8jl3bXqKxr1iYurIKttrxTl+32psabHaYtHhlymZpxrDivwOJLKd282kNF2h
+wV7Yl3V5QHw3960GyF+J7K0s/Kp4mKFmtnpNhfwbKwwkULkKmiS0iVllpqFLqE+P0fsIP5Eaeth
4aNS+Eehkb7lpVGevI4Qi327JnwnwS6G/DZSUVU7
`protect end_protected
